`timescale 1 ns/1 ps
`include "SRAM_SP_ADV.v"

module hw4(CLK, WA, A_CPU, WorC, CEN, D, Hit, Q);

input CLK;
input [5:0]WA;
input [15:0]A_CPU;
input WorC;
input CEN;
input [127:0]D;
output wire Hit;
output wire [127:0]Q;

reg [2:0]EMA=3'b000;

reg [7:0]A;

reg [15:0]CAM[63:0];
reg [63:0]valid;

wire [5:0]encoder;

always @(posedge CLK)begin
    case(WA)
    6'b000000:begin
    if(~WorC)
        CAM[0][15:0]<=A_CPU[15:0];
    else
        CAM[0][15:0]<=CAM[0][15:0];
    end
    6'b000001:begin
    if(~WorC)
        CAM[1][15:0]<=A_CPU[15:0];
    else
        CAM[1][15:0]<=CAM[1][15:0];
    end
    6'b000010:begin
    if(~WorC)
        CAM[2][15:0]<=A_CPU[15:0];
    else
        CAM[2][15:0]<=CAM[2][15:0];
    end
    6'b000011:begin
    if(~WorC)
        CAM[3][15:0]<=A_CPU[15:0];
    else
        CAM[3][15:0]<=CAM[3][15:0];
    end
    6'b000100:begin
    if(~WorC)
        CAM[4][15:0]<=A_CPU[15:0];
    else
        CAM[4][15:0]<=CAM[4][15:0];
    end
    6'b000101:begin
    if(~WorC)
        CAM[5][15:0]<=A_CPU[15:0];
    else
        CAM[5][15:0]<=CAM[5][15:0];
    end
    6'b000110:begin
    if(~WorC)
        CAM[6][15:0]<=A_CPU[15:0];
    else
        CAM[6][15:0]<=CAM[6][15:0];
    end
    6'b000111:begin
    if(~WorC)
        CAM[7][15:0]<=A_CPU[15:0];
    else
        CAM[7][15:0]<=CAM[7][15:0];
    end
    6'b001000:begin
    if(~WorC)
        CAM[8][15:0]<=A_CPU[15:0];
    else
        CAM[8][15:0]<=CAM[8][15:0];
    end
    6'b001001:begin
    if(~WorC)
        CAM[9][15:0]<=A_CPU[15:0];
    else
        CAM[9][15:0]<=CAM[9][15:0];
    end
    6'b001010:begin
    if(~WorC)
        CAM[10][15:0]<=A_CPU[15:0];
    else
        CAM[10][15:0]<=CAM[10][15:0];
    end
    6'b001011:begin
    if(~WorC)
        CAM[11][15:0]<=A_CPU[15:0];
    else
        CAM[11][15:0]<=CAM[11][15:0];
    end
    6'b001100:begin
    if(~WorC)
        CAM[12][15:0]<=A_CPU[15:0];
    else
        CAM[12][15:0]<=CAM[12][15:0];
    end
    6'b001101:begin
    if(~WorC)
        CAM[13][15:0]<=A_CPU[15:0];
    else
        CAM[13][15:0]<=CAM[13][15:0];
    end
    6'b001110:begin
    if(~WorC)
        CAM[14][15:0]<=A_CPU[15:0];
    else
        CAM[14][15:0]<=CAM[14][15:0];
    end
    6'b001111:begin
    if(~WorC)
        CAM[15][15:0]<=A_CPU[15:0];
    else
        CAM[15][15:0]<=CAM[15][15:0];
    end
    6'b010000:begin
    if(~WorC)
        CAM[16][15:0]<=A_CPU[15:0];
    else
        CAM[16][15:0]<=CAM[16][15:0];
    end
    6'b010001:begin
    if(~WorC)
        CAM[17][15:0]<=A_CPU[15:0];
    else
        CAM[17][15:0]<=CAM[17][15:0];
    end
    6'b010010:begin
    if(~WorC)
        CAM[18][15:0]<=A_CPU[15:0];
    else
        CAM[18][15:0]<=CAM[18][15:0];
    end
    6'b010011:begin
    if(~WorC)
        CAM[19][15:0]<=A_CPU[15:0];
    else
        CAM[19][15:0]<=CAM[19][15:0];
    end
    6'b010100:begin
    if(~WorC)
        CAM[20][15:0]<=A_CPU[15:0];
    else
        CAM[20][15:0]<=CAM[20][15:0];
    end
    6'b010101:begin
    if(~WorC)
        CAM[21][15:0]<=A_CPU[15:0];
    else
        CAM[21][15:0]<=CAM[21][15:0];
    end
    6'b010110:begin
    if(~WorC)
        CAM[22][15:0]<=A_CPU[15:0];
    else
        CAM[22][15:0]<=CAM[22][15:0];
    end
    6'b010111:begin
    if(~WorC)
        CAM[23][15:0]<=A_CPU[15:0];
    else
        CAM[23][15:0]<=CAM[23][15:0];
    end
    6'b011000:begin
    if(~WorC)
        CAM[24][15:0]<=A_CPU[15:0];
    else
        CAM[24][15:0]<=CAM[24][15:0];
    end
    6'b011001:begin
    if(~WorC)
        CAM[25][15:0]<=A_CPU[15:0];
    else
        CAM[25][15:0]<=CAM[25][15:0];
    end
    6'b011010:begin
    if(~WorC)
        CAM[26][15:0]<=A_CPU[15:0];
    else
        CAM[26][15:0]<=CAM[26][15:0];
    end
    6'b011011:begin
    if(~WorC)
        CAM[27][15:0]<=A_CPU[15:0];
    else
        CAM[27][15:0]<=CAM[27][15:0];
    end
    6'b011100:begin
    if(~WorC)
        CAM[28][15:0]<=A_CPU[15:0];
    else
        CAM[28][15:0]<=CAM[28][15:0];
    end
    6'b011101:begin
    if(~WorC)
        CAM[29][15:0]<=A_CPU[15:0];
    else
        CAM[29][15:0]<=CAM[29][15:0];
    end
    6'b011110:begin
    if(~WorC)
        CAM[30][15:0]<=A_CPU[15:0];
    else
        CAM[30][15:0]<=CAM[30][15:0];
    end
    6'b011111:begin
    if(~WorC)
        CAM[31][15:0]<=A_CPU[15:0];
    else
        CAM[31][15:0]<=CAM[31][15:0];
    end
    6'b100000:begin
    if(~WorC)
        CAM[32][15:0]<=A_CPU[15:0];
    else
        CAM[32][15:0]<=CAM[32][15:0];
    end
    6'b100001:begin
    if(~WorC)
        CAM[33][15:0]<=A_CPU[15:0];
    else
        CAM[33][15:0]<=CAM[33][15:0];
    end
    6'b100010:begin
    if(~WorC)
        CAM[34][15:0]<=A_CPU[15:0];
    else
        CAM[34][15:0]<=CAM[34][15:0];
    end
    6'b100011:begin
    if(~WorC)
        CAM[35][15:0]<=A_CPU[15:0];
    else
        CAM[35][15:0]<=CAM[35][15:0];
    end
    6'b100100:begin
    if(~WorC)
        CAM[36][15:0]<=A_CPU[15:0];
    else
        CAM[36][15:0]<=CAM[36][15:0];
    end
    6'b100101:begin
    if(~WorC)
        CAM[37][15:0]<=A_CPU[15:0];
    else
        CAM[37][15:0]<=CAM[37][15:0];
    end
    6'b100110:begin
    if(~WorC)
        CAM[38][15:0]<=A_CPU[15:0];
    else
        CAM[38][15:0]<=CAM[38][15:0];
    end
    6'b100111:begin
    if(~WorC)
        CAM[39][15:0]<=A_CPU[15:0];
    else
        CAM[39][15:0]<=CAM[39][15:0];
    end
    6'b101000:begin
    if(~WorC)
        CAM[40][15:0]<=A_CPU[15:0];
    else
        CAM[40][15:0]<=CAM[40][15:0];
    end
    6'b101001:begin
    if(~WorC)
        CAM[41][15:0]<=A_CPU[15:0];
    else
        CAM[41][15:0]<=CAM[41][15:0];
    end
    6'b101010:begin
    if(~WorC)
        CAM[42][15:0]<=A_CPU[15:0];
    else
        CAM[42][15:0]<=CAM[42][15:0];
    end
    6'b101011:begin
    if(~WorC)
        CAM[43][15:0]<=A_CPU[15:0];
    else
        CAM[43][15:0]<=CAM[43][15:0];
    end
    6'b101100:begin
    if(~WorC)
        CAM[44][15:0]<=A_CPU[15:0];
    else
        CAM[44][15:0]<=CAM[44][15:0];
    end
    6'b101101:begin
    if(~WorC)
        CAM[45][15:0]<=A_CPU[15:0];
    else
        CAM[45][15:0]<=CAM[45][15:0];
    end
    6'b101110:begin
    if(~WorC)
        CAM[46][15:0]<=A_CPU[15:0];
    else
        CAM[46][15:0]<=CAM[46][15:0];
    end
    6'b101111:begin
    if(~WorC)
        CAM[47][15:0]<=A_CPU[15:0];
    else
        CAM[47][15:0]<=CAM[47][15:0];
    end
    6'b110000:begin
    if(~WorC)
        CAM[48][15:0]<=A_CPU[15:0];
    else
        CAM[48][15:0]<=CAM[48][15:0];
    end
    6'b110001:begin
    if(~WorC)
        CAM[49][15:0]<=A_CPU[15:0];
    else
        CAM[49][15:0]<=CAM[49][15:0];
    end
    6'b110010:begin
    if(~WorC)
        CAM[50][15:0]<=A_CPU[15:0];
    else
        CAM[50][15:0]<=CAM[50][15:0];
    end
    6'b110011:begin
    if(~WorC)
        CAM[51][15:0]<=A_CPU[15:0];
    else
        CAM[51][15:0]<=CAM[51][15:0];
    end
    6'b110100:begin
    if(~WorC)
        CAM[52][15:0]<=A_CPU[15:0];
    else
        CAM[52][15:0]<=CAM[52][15:0];
    end
    6'b110101:begin
    if(~WorC)
        CAM[53][15:0]<=A_CPU[15:0];
    else
        CAM[53][15:0]<=CAM[53][15:0];
    end
    6'b110110:begin
    if(~WorC)
        CAM[54][15:0]<=A_CPU[15:0];
    else
        CAM[54][15:0]<=CAM[54][15:0];
    end
    6'b110111:begin
    if(~WorC)
        CAM[55][15:0]<=A_CPU[15:0];
    else
        CAM[55][15:0]<=CAM[55][15:0];
    end
    6'b111000:begin
    if(~WorC)
        CAM[56][15:0]<=A_CPU[15:0];
    else
        CAM[56][15:0]<=CAM[56][15:0];
    end
    6'b111001:begin
    if(~WorC)
        CAM[57][15:0]<=A_CPU[15:0];
    else
        CAM[57][15:0]<=CAM[57][15:0];
    end
    6'b111010:begin
    if(~WorC)
        CAM[58][15:0]<=A_CPU[15:0];
    else
        CAM[58][15:0]<=CAM[58][15:0];
    end
    6'b111011:begin
    if(~WorC)
        CAM[59][15:0]<=A_CPU[15:0];
    else
        CAM[59][15:0]<=CAM[59][15:0];
    end
    6'b111100:begin
    if(~WorC)
        CAM[60][15:0]<=A_CPU[15:0];
    else
        CAM[60][15:0]<=CAM[60][15:0];
    end
    6'b111101:begin
    if(~WorC)
        CAM[61][15:0]<=A_CPU[15:0];
    else
        CAM[61][15:0]<=CAM[61][15:0];
    end
    6'b111110:begin
    if(~WorC)
        CAM[62][15:0]<=A_CPU[15:0];
    else
        CAM[62][15:0]<=CAM[62][15:0];
    end
    6'b111111:begin
    if(~WorC)
        CAM[63][15:0]<=A_CPU[15:0];
    else
        CAM[63][15:0]<=CAM[63][15:0];
    end
    endcase
end

always @(WorC, A_CPU)begin
    case(A_CPU)
    CAM[0][15:0]:
    if(WorC)begin
        valid[63:1]=1'b0;
        valid[0]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[1][15:0]:
    if(WorC)begin
        valid[0]=1'b0;
        valid[63:2]=1'b0;
        valid[1]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[2][15:0]:
    if(WorC)begin
        valid[1:0]=1'b0;
        valid[63:3]=1'b0;
        valid[2]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[3][15:0]:
    if(WorC)begin
        valid[2:0]=1'b0;
        valid[63:4]=1'b0;
        valid[3]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[4][15:0]:
    if(WorC)begin
        valid[3:0]=1'b0;
        valid[63:5]=1'b0;
        valid[4]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[5][15:0]:
    if(WorC)begin
        valid[4:0]=1'b0;
        valid[63:6]=1'b0;
        valid[5]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[6][15:0]:
    if(WorC)begin
        valid[5:0]=1'b0;
        valid[63:7]=1'b0;
        valid[6]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[7][15:0]:
    if(WorC)begin
        valid[6:0]=1'b0;
        valid[63:8]=1'b0;
        valid[7]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[8][15:0]:
    if(WorC)begin
        valid[7:0]=1'b0;
        valid[63:9]=1'b0;
        valid[8]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[9][15:0]:
    if(WorC)begin
        valid[8:0]=1'b0;
        valid[63:10]=1'b0;
        valid[9]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[10][15:0]:
    if(WorC)begin
        valid[9:0]=1'b0;
        valid[63:11]=1'b0;
        valid[10]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[11][15:0]:
    if(WorC)begin
        valid[10:0]=1'b0;
        valid[63:12]=1'b0;
        valid[11]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[12][15:0]:
    if(WorC)begin
        valid[11:0]=1'b0;
        valid[63:13]=1'b0;
        valid[12]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[13][15:0]:
    if(WorC)begin
        valid[12:0]=1'b0;
        valid[63:14]=1'b0;
        valid[13]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[14][15:0]:
    if(WorC)begin
        valid[13:0]=1'b0;
        valid[63:15]=1'b0;
        valid[14]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[15][15:0]:
    if(WorC)begin
        valid[14:0]=1'b0;
        valid[63:16]=1'b0;
        valid[15]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[16][15:0]:
    if(WorC)begin
        valid[15:0]=1'b0;
        valid[63:17]=1'b0;
        valid[16]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[17][15:0]:
    if(WorC)begin
        valid[16:0]=1'b0;
        valid[63:18]=1'b0;
        valid[17]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[18][15:0]:
    if(WorC)begin
        valid[17:0]=1'b0;
        valid[63:19]=1'b0;
        valid[18]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[19][15:0]:
    if(WorC)begin
        valid[18:0]=1'b0;
        valid[63:20]=1'b0;
        valid[19]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[20][15:0]:
    if(WorC)begin
        valid[19:0]=1'b0;
        valid[63:21]=1'b0;
        valid[20]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[21][15:0]:
    if(WorC)begin
        valid[20:0]=1'b0;
        valid[63:22]=1'b0;
        valid[21]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[22][15:0]:
    if(WorC)begin
        valid[21:0]=1'b0;
        valid[63:23]=1'b0;
        valid[22]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[23][15:0]:
    if(WorC)begin
        valid[22:0]=1'b0;
        valid[63:24]=1'b0;
        valid[23]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[24][15:0]:
    if(WorC)begin
        valid[23:0]=1'b0;
        valid[63:25]=1'b0;
        valid[24]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[25][15:0]:
    if(WorC)begin
        valid[24:0]=1'b0;
        valid[63:26]=1'b0;
        valid[25]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[26][15:0]:
    if(WorC)begin
        valid[25:0]=1'b0;
        valid[63:27]=1'b0;
        valid[26]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[27][15:0]:
    if(WorC)begin
        valid[26:0]=1'b0;
        valid[63:28]=1'b0;
        valid[27]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[28][15:0]:
    if(WorC)begin
        valid[27:0]=1'b0;
        valid[63:29]=1'b0;
        valid[28]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[29][15:0]:
    if(WorC)begin
        valid[28:0]=1'b0;
        valid[63:30]=1'b0;
        valid[29]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[30][15:0]:
    if(WorC)begin
        valid[29:0]=1'b0;
        valid[63:31]=1'b0;
        valid[30]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[31][15:0]:
    if(WorC)begin
        valid[30:0]=1'b0;
        valid[63:32]=1'b0;
        valid[31]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[32][15:0]:
    if(WorC)begin
        valid[31:0]=1'b0;
        valid[63:33]=1'b0;
        valid[32]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[33][15:0]:
    if(WorC)begin
        valid[32:0]=1'b0;
        valid[63:34]=1'b0;
        valid[33]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[34][15:0]:
    if(WorC)begin
        valid[33:0]=1'b0;
        valid[63:35]=1'b0;
        valid[34]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[35][15:0]:
    if(WorC)begin
        valid[34:0]=1'b0;
        valid[63:36]=1'b0;
        valid[35]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[36][15:0]:
    if(WorC)begin
        valid[35:0]=1'b0;
        valid[63:37]=1'b0;
        valid[36]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[37][15:0]:
    if(WorC)begin
        valid[36:0]=1'b0;
        valid[63:38]=1'b0;
        valid[37]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[38][15:0]:
    if(WorC)begin
        valid[37:0]=1'b0;
        valid[63:39]=1'b0;
        valid[38]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[39][15:0]:
    if(WorC)begin
        valid[38:0]=1'b0;
        valid[63:40]=1'b0;
        valid[39]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[40][15:0]:
    if(WorC)begin
        valid[39:0]=1'b0;
        valid[63:41]=1'b0;
        valid[40]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[41][15:0]:
    if(WorC)begin
        valid[40:0]=1'b0;
        valid[63:42]=1'b0;
        valid[41]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[42][15:0]:
    if(WorC)begin
        valid[41:0]=1'b0;
        valid[63:43]=1'b0;
        valid[42]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[43][15:0]:
    if(WorC)begin
        valid[42:0]=1'b0;
        valid[63:44]=1'b0;
        valid[43]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[44][15:0]:
    if(WorC)begin
        valid[43:0]=1'b0;
        valid[63:45]=1'b0;
        valid[44]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[45][15:0]:
    if(WorC)begin
        valid[44:0]=1'b0;
        valid[63:46]=1'b0;
        valid[45]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[46][15:0]:
    if(WorC)begin
        valid[45:0]=1'b0;
        valid[63:47]=1'b0;
        valid[46]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[47][15:0]:
    if(WorC)begin
        valid[46:0]=1'b0;
        valid[63:48]=1'b0;
        valid[47]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[48][15:0]:
    if(WorC)begin
        valid[47:0]=1'b0;
        valid[63:49]=1'b0;
        valid[48]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[49][15:0]:
    if(WorC)begin
        valid[48:0]=1'b0;
        valid[63:50]=1'b0;
        valid[49]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[50][15:0]:
    if(WorC)begin
        valid[49:0]=1'b0;
        valid[63:51]=1'b0;
        valid[50]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[51][15:0]:
    if(WorC)begin
        valid[50:0]=1'b0;
        valid[63:52]=1'b0;
        valid[51]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[52][15:0]:
    if(WorC)begin
        valid[51:0]=1'b0;
        valid[63:53]=1'b0;
        valid[52]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[53][15:0]:
    if(WorC)begin
        valid[52:0]=1'b0;
        valid[63:54]=1'b0;
        valid[53]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[54][15:0]:
    if(WorC)begin
        valid[53:0]=1'b0;
        valid[63:55]=1'b0;
        valid[54]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[55][15:0]:
    if(WorC)begin
        valid[54:0]=1'b0;
        valid[63:56]=1'b0;
        valid[55]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[56][15:0]:
    if(WorC)begin
        valid[55:0]=1'b0;
        valid[63:57]=1'b0;
        valid[56]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[57][15:0]:
    if(WorC)begin
        valid[56:0]=1'b0;
        valid[63:58]=1'b0;
        valid[57]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[58][15:0]:
    if(WorC)begin
        valid[57:0]=1'b0;
        valid[63:59]=1'b0;
        valid[58]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[59][15:0]:
    if(WorC)begin
        valid[58:0]=1'b0;
        valid[63:60]=1'b0;
        valid[59]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[60][15:0]:
    if(WorC)begin
        valid[59:0]=1'b0;
        valid[63:61]=1'b0;
        valid[60]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[61][15:0]:
    if(WorC)begin
        valid[60:0]=1'b0;
        valid[63:62]=1'b0;
        valid[61]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[62][15:0]:
    if(WorC)begin
        valid[61:0]=1'b0;
        valid[63]=1'b0;
        valid[62]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    CAM[63][15:0]:
    if(WorC)begin
        valid[62:0]=1'b0;
        valid[63]=1'b1;
    end
    else
        valid[63:0]=64'b0;
    default:valid[63:0]=64'b0;
    endcase
end

assign Hit=(|valid);

assign encoder[0]=valid[1]||valid[3]||valid[5]||valid[7]||valid[9]||valid[11]||valid[13]||valid[15]||valid[17]||valid[19]||valid[21]||valid[23]||valid[25]||valid[27]||valid[29]||valid[31]||valid[33]||valid[35]||valid[37]||valid[39]||valid[41]||valid[43]||valid[45]||valid[47]||valid[49]||valid[51]||valid[53]||valid[55]||valid[57]||valid[59]||valid[61]||valid[63];
assign encoder[1]=valid[2]||valid[3]||valid[6]||valid[7]||valid[10]||valid[11]||valid[14]||valid[15]||valid[18]||valid[19]||valid[22]||valid[23]||valid[26]||valid[27]||valid[30]||valid[31]||valid[34]||valid[35]||valid[38]||valid[39]||valid[42]||valid[43]||valid[46]||valid[47]||valid[50]||valid[51]||valid[54]||valid[55]||valid[58]||valid[59]||valid[62]||valid[63];
assign encoder[2]=valid[4]||valid[5]||valid[6]||valid[7]||valid[12]||valid[13]||valid[14]||valid[15]||valid[20]||valid[21]||valid[22]||valid[23]||valid[28]||valid[29]||valid[30]||valid[31]||valid[36]||valid[37]||valid[38]||valid[39]||valid[44]||valid[45]||valid[46]||valid[47]||valid[52]||valid[53]||valid[54]||valid[55]||valid[60]||valid[61]||valid[62]||valid[63];
assign encoder[3]=valid[8]||valid[9]||valid[10]||valid[11]||valid[12]||valid[13]||valid[14]||valid[15]||valid[24]||valid[25]||valid[26]||valid[27]||valid[28]||valid[29]||valid[30]||valid[31]||valid[40]||valid[41]||valid[42]||valid[43]||valid[44]||valid[45]||valid[46]||valid[47]||valid[56]||valid[57]||valid[58]||valid[59]||valid[60]||valid[61]||valid[62]||valid[63];
assign encoder[4]=valid[16]||valid[17]||valid[18]||valid[19]||valid[20]||valid[21]||valid[22]||valid[23]||valid[24]||valid[25]||valid[26]||valid[27]||valid[28]||valid[29]||valid[30]||valid[31]||valid[48]||valid[49]||valid[50]||valid[51]||valid[52]||valid[53]||valid[54]||valid[55]||valid[56]||valid[57]||valid[58]||valid[59]||valid[60]||valid[61]||valid[62]||valid[63];
assign encoder[5]=(|valid[63:32]);



always @(valid, WorC, WA, encoder)begin
    if(~WorC)
        A[7:0]={2'b0, WA};
    else if(|valid)
        A[7:0]={2'b0, encoder};
    else
        A[7:0]=8'b11111111;
end

SRAM_SP_ADV S0(.Q(Q), .CLK(~CLK), .CEN(CEN), .WEN(WorC), .A(A), .D(D), .EMA(EMA));

endmodule