.SUBCKT DCIM VSS VDD clk rst_n in_valid in_data1[127] in_data1[126] in_data1[125] in_data1[124] in_data1[123] in_data1[122] in_data1[121] in_data1[120] in_data1[119] in_data1[118] in_data1[117] in_data1[116] in_data1[115] in_data1[114] in_data1[113] in_data1[112] in_data1[111] in_data1[110] in_data1[109] in_data1[108] in_data1[107] in_data1[106] in_data1[105] in_data1[104] in_data1[103] in_data1[102] in_data1[101] in_data1[100] in_data1[99] in_data1[98] in_data1[97] in_data1[96] in_data1[95] in_data1[94] in_data1[93] in_data1[92] in_data1[91] in_data1[90] in_data1[89] in_data1[88] in_data1[87] in_data1[86] in_data1[85] in_data1[84] in_data1[83] in_data1[82] in_data1[81] in_data1[80] in_data1[79] in_data1[78] in_data1[77] in_data1[76] in_data1[75] in_data1[74] in_data1[73] in_data1[72] in_data1[71] in_data1[70] in_data1[69] in_data1[68] in_data1[67] in_data1[66] in_data1[65] in_data1[64] in_data1[63] in_data1[62] in_data1[61] in_data1[60] in_data1[59] in_data1[58] in_data1[57] in_data1[56] in_data1[55] in_data1[54] in_data1[53] in_data1[52] in_data1[51] in_data1[50] in_data1[49] in_data1[48] in_data1[47] in_data1[46] in_data1[45] in_data1[44] in_data1[43] in_data1[42] in_data1[41] in_data1[40] in_data1[39] in_data1[38] in_data1[37] in_data1[36] in_data1[35] in_data1[34] in_data1[33] in_data1[32] in_data1[31] in_data1[30] in_data1[29] in_data1[28] in_data1[27] in_data1[26] in_data1[25] in_data1[24] in_data1[23] in_data1[22] in_data1[21] in_data1[20] in_data1[19] in_data1[18] in_data1[17] in_data1[16] in_data1[15] in_data1[14] in_data1[13] in_data1[12] in_data1[11] in_data1[10] in_data1[9] in_data1[8] in_data1[7] in_data1[6] in_data1[5] in_data1[4] in_data1[3] in_data1[2] in_data1[1] in_data1[0] in_data2[127] in_data2[126] in_data2[125] in_data2[124] in_data2[123] in_data2[122] in_data2[121] in_data2[120] in_data2[119] in_data2[118] in_data2[117] in_data2[116] in_data2[115] in_data2[114] in_data2[113] in_data2[112] in_data2[111] in_data2[110] in_data2[109] in_data2[108] in_data2[107] in_data2[106] in_data2[105] in_data2[104] in_data2[103] in_data2[102] in_data2[101] in_data2[100] in_data2[99] in_data2[98] in_data2[97] in_data2[96] in_data2[95] in_data2[94] in_data2[93] in_data2[92] in_data2[91] in_data2[90] in_data2[89] in_data2[88] in_data2[87] in_data2[86] in_data2[85] in_data2[84] in_data2[83] in_data2[82] in_data2[81] in_data2[80] in_data2[79] in_data2[78] in_data2[77] in_data2[76] in_data2[75] in_data2[74] in_data2[73] in_data2[72] in_data2[71] in_data2[70] in_data2[69] in_data2[68] in_data2[67] in_data2[66] in_data2[65] in_data2[64] in_data2[63] in_data2[62] in_data2[61] in_data2[60] in_data2[59] in_data2[58] in_data2[57] in_data2[56] in_data2[55] in_data2[54] in_data2[53] in_data2[52] in_data2[51] in_data2[50] in_data2[49] in_data2[48] in_data2[47] in_data2[46] in_data2[45] in_data2[44] in_data2[43] in_data2[42] in_data2[41] in_data2[40] in_data2[39] in_data2[38] in_data2[37] in_data2[36] in_data2[35] in_data2[34] in_data2[33] in_data2[32] in_data2[31] in_data2[30] in_data2[29] in_data2[28] in_data2[27] in_data2[26] in_data2[25] in_data2[24] in_data2[23] in_data2[22] in_data2[21] in_data2[20] in_data2[19] in_data2[18] in_data2[17] in_data2[16] in_data2[15] in_data2[14] in_data2[13] in_data2[12] in_data2[11] in_data2[10] in_data2[9] in_data2[8] in_data2[7] in_data2[6] in_data2[5] in_data2[4] in_data2[3] in_data2[2] in_data2[1] in_data2[0] in_data3[127] in_data3[126] in_data3[125] in_data3[124] in_data3[123] in_data3[122] in_data3[121] in_data3[120] in_data3[119] in_data3[118] in_data3[117] in_data3[116] in_data3[115] in_data3[114] in_data3[113] in_data3[112] in_data3[111] in_data3[110] in_data3[109] in_data3[108] in_data3[107] in_data3[106] in_data3[105] in_data3[104] in_data3[103] in_data3[102] in_data3[101] in_data3[100] in_data3[99] in_data3[98] in_data3[97] in_data3[96] in_data3[95] in_data3[94] in_data3[93] in_data3[92] in_data3[91] in_data3[90] in_data3[89] in_data3[88] in_data3[87] in_data3[86] in_data3[85] in_data3[84] in_data3[83] in_data3[82] in_data3[81] in_data3[80] in_data3[79] in_data3[78] in_data3[77] in_data3[76] in_data3[75] in_data3[74] in_data3[73] in_data3[72] in_data3[71] in_data3[70] in_data3[69] in_data3[68] in_data3[67] in_data3[66] in_data3[65] in_data3[64] in_data3[63] in_data3[62] in_data3[61] in_data3[60] in_data3[59] in_data3[58] in_data3[57] in_data3[56] in_data3[55] in_data3[54] in_data3[53] in_data3[52] in_data3[51] in_data3[50] in_data3[49] in_data3[48] in_data3[47] in_data3[46] in_data3[45] in_data3[44] in_data3[43] in_data3[42] in_data3[41] in_data3[40] in_data3[39] in_data3[38] in_data3[37] in_data3[36] in_data3[35] in_data3[34] in_data3[33] in_data3[32] in_data3[31] in_data3[30] in_data3[29] in_data3[28] in_data3[27] in_data3[26] in_data3[25] in_data3[24] in_data3[23] in_data3[22] in_data3[21] in_data3[20] in_data3[19] in_data3[18] in_data3[17] in_data3[16] in_data3[15] in_data3[14] in_data3[13] in_data3[12] in_data3[11] in_data3[10] in_data3[9] in_data3[8] in_data3[7] in_data3[6] in_data3[5] in_data3[4] in_data3[3] in_data3[2] in_data3[1] in_data3[0] in_data4[127] in_data4[126] in_data4[125] in_data4[124] in_data4[123] in_data4[122] in_data4[121] in_data4[120] in_data4[119] in_data4[118] in_data4[117] in_data4[116] in_data4[115] in_data4[114] in_data4[113] in_data4[112] in_data4[111] in_data4[110] in_data4[109] in_data4[108] in_data4[107] in_data4[106] in_data4[105] in_data4[104] in_data4[103] in_data4[102] in_data4[101] in_data4[100] in_data4[99] in_data4[98] in_data4[97] in_data4[96] in_data4[95] in_data4[94] in_data4[93] in_data4[92] in_data4[91] in_data4[90] in_data4[89] in_data4[88] in_data4[87] in_data4[86] in_data4[85] in_data4[84] in_data4[83] in_data4[82] in_data4[81] in_data4[80] in_data4[79] in_data4[78] in_data4[77] in_data4[76] in_data4[75] in_data4[74] in_data4[73] in_data4[72] in_data4[71] in_data4[70] in_data4[69] in_data4[68] in_data4[67] in_data4[66] in_data4[65] in_data4[64] in_data4[63] in_data4[62] in_data4[61] in_data4[60] in_data4[59] in_data4[58] in_data4[57] in_data4[56] in_data4[55] in_data4[54] in_data4[53] in_data4[52] in_data4[51] in_data4[50] in_data4[49] in_data4[48] in_data4[47] in_data4[46] in_data4[45] in_data4[44] in_data4[43] in_data4[42] in_data4[41] in_data4[40] in_data4[39] in_data4[38] in_data4[37] in_data4[36] in_data4[35] in_data4[34] in_data4[33] in_data4[32] in_data4[31] in_data4[30] in_data4[29] in_data4[28] in_data4[27] in_data4[26] in_data4[25] in_data4[24] in_data4[23] in_data4[22] in_data4[21] in_data4[20] in_data4[19] in_data4[18] in_data4[17] in_data4[16] in_data4[15] in_data4[14] in_data4[13] in_data4[12] in_data4[11] in_data4[10] in_data4[9] in_data4[8] in_data4[7] in_data4[6] in_data4[5] in_data4[4] in_data4[3] in_data4[2] in_data4[1] in_data4[0] out_valid O1[12] O1[11] O1[10] O1[9] O1[8] O1[7] O1[6] O1[5] O1[4] O1[3] O1[2] O1[1] O1[0] O2[12] O2[11] O2[10] O2[9] O2[8] O2[7] O2[6] O2[5] O2[4] O2[3] O2[2] O2[1] O2[0] O3[12] O3[11] O3[10] O3[9] O3[8] O3[7] O3[6] O3[5] O3[4] O3[3] O3[2] O3[1] O3[0] O4[12] O4[11] O4[10] O4[9] O4[8] O4[7] O4[6] O4[5] O4[4] O4[3] O4[2] O4[1] O4[0]
XU1157 VSS VDD n287 n289 n1074 AND2x2_ASAP7_75t_R
Xin_valid_dff_reg VSS VDD clk in_valid n183 n938 n345 ASYNC_DFFHx1_ASAP7_75t_R
Xin_valid_dff_2_reg VSS VDD clk n860 n183 n872 n344 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_12_ VSS VDD clk N1614 n183 n870 n343 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_11_ VSS VDD clk N1613 n183 n944 n342 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_10_ VSS VDD clk N1612 n183 n890 n341 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_9_ VSS VDD clk N1611 n183 n918 n340 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_8_ VSS VDD clk N1610 n183 n902 n339 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_7_ VSS VDD clk N1609 n183 n952 n338 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_6_ VSS VDD clk N1608 n183 n876 n337 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_5_ VSS VDD clk N1607 n183 n978 n336 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_4_ VSS VDD clk N1606 n183 n1015 n335 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_3_ VSS VDD clk N1605 n183 n949 n334 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_2_ VSS VDD clk N1604 n183 n931 n333 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_1_ VSS VDD clk N1603 n183 n979 n332 ASYNC_DFFHx1_ASAP7_75t_R
XO4_reg_0_ VSS VDD clk N1602 n183 n959 n331 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_12_ VSS VDD clk N1575 n183 n885 n330 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_11_ VSS VDD clk N1574 n183 n903 n329 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_10_ VSS VDD clk N1573 n183 n905 n328 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_9_ VSS VDD clk N1572 n183 n958 n327 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_8_ VSS VDD clk N1571 n183 n981 n326 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_7_ VSS VDD clk N1570 n183 n986 n325 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_6_ VSS VDD clk N1569 n183 n988 n324 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_5_ VSS VDD clk N1568 n183 n875 n323 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_4_ VSS VDD clk N1567 n183 n940 n322 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_3_ VSS VDD clk N1566 n183 n881 n321 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_2_ VSS VDD clk N1565 n183 n873 n320 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_1_ VSS VDD clk N1564 n183 n866 n319 ASYNC_DFFHx1_ASAP7_75t_R
XO1_reg_0_ VSS VDD clk N1563 n183 n927 n318 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_12_ VSS VDD clk N1588 n183 n972 n317 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_11_ VSS VDD clk N1587 n183 n867 n316 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_10_ VSS VDD clk N1586 n183 n884 n315 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_9_ VSS VDD clk N1585 n183 n1007 n314 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_8_ VSS VDD clk N1584 n183 n982 n313 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_7_ VSS VDD clk N1583 n183 n976 n312 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_6_ VSS VDD clk N1582 n183 n962 n311 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_5_ VSS VDD clk N1581 n183 n898 n310 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_4_ VSS VDD clk N1580 n183 n985 n309 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_3_ VSS VDD clk N1579 n183 n871 n308 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_2_ VSS VDD clk N1578 n183 n864 n307 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_1_ VSS VDD clk N1577 n183 n874 n306 ASYNC_DFFHx1_ASAP7_75t_R
XO2_reg_0_ VSS VDD clk N1576 n183 n920 n305 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_12_ VSS VDD clk N1601 n183 n951 n304 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_11_ VSS VDD clk N1600 n183 n939 n303 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_10_ VSS VDD clk N1599 n183 n891 n302 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_9_ VSS VDD clk N1598 n183 n987 n301 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_8_ VSS VDD clk N1597 n183 n921 n300 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_7_ VSS VDD clk N1596 n183 n908 n299 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_6_ VSS VDD clk N1595 n183 n897 n298 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_5_ VSS VDD clk N1594 n183 n877 n297 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_4_ VSS VDD clk N1593 n183 n880 n296 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_3_ VSS VDD clk N1592 n183 n923 n295 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_2_ VSS VDD clk N1591 n183 n879 n294 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_1_ VSS VDD clk N1590 n183 n889 n293 ASYNC_DFFHx1_ASAP7_75t_R
XO3_reg_0_ VSS VDD clk N1589 n183 n1008 n292 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg VSS VDD clk n863 n183 n932 n291 ASYNC_DFFHx1_ASAP7_75t_R
Xcnt_reg_0_ VSS VDD clk n290 n183 n865 n289 ASYNC_DFFHx1_ASAP7_75t_R
Xcnt_reg_1_ VSS VDD clk n288 n183 n1012 n287 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_12_ VSS VDD clk n286 n183 n983 n285 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_11_ VSS VDD clk n284 n183 n930 n283 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_10_ VSS VDD clk n282 n183 n893 n281 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_9_ VSS VDD clk n280 n183 n909 n279 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_8_ VSS VDD clk n278 n183 n1001 n277 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_7_ VSS VDD clk n276 n183 n953 n275 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_6_ VSS VDD clk n274 n183 n892 n273 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_5_ VSS VDD clk n272 n183 n906 n271 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_4_ VSS VDD clk n270 n183 n894 n269 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_3_ VSS VDD clk n268 n183 n1018 n267 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_2_ VSS VDD clk n266 n183 n954 n265 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_1_ VSS VDD clk n264 n183 n977 n263 ASYNC_DFFHx1_ASAP7_75t_R
Xsum4_reg_0_ VSS VDD clk n262 n183 n945 n261 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_12_ VSS VDD clk n260 n183 n904 n259 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_11_ VSS VDD clk n258 n183 n896 n257 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_10_ VSS VDD clk n256 n183 n947 n255 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_9_ VSS VDD clk n254 n183 n887 n253 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_8_ VSS VDD clk n252 n183 n899 n251 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_7_ VSS VDD clk n250 n183 n1013 n249 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_6_ VSS VDD clk n248 n183 n924 n247 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_5_ VSS VDD clk n246 n183 n878 n245 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_4_ VSS VDD clk n244 n183 n1006 n243 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_3_ VSS VDD clk n242 n183 n922 n241 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_2_ VSS VDD clk n240 n183 n963 n239 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_1_ VSS VDD clk n238 n183 n895 n237 ASYNC_DFFHx1_ASAP7_75t_R
Xsum1_reg_0_ VSS VDD clk n236 n183 n950 n235 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_12_ VSS VDD clk n234 n183 n1014 n233 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_11_ VSS VDD clk n232 n183 n1011 n231 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_10_ VSS VDD clk n230 n183 n948 n229 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_9_ VSS VDD clk n228 n183 n973 n227 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_8_ VSS VDD clk n226 n183 n942 n225 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_7_ VSS VDD clk n224 n183 n1010 n223 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_6_ VSS VDD clk n222 n183 n925 n221 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_5_ VSS VDD clk n220 n183 n869 n219 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_4_ VSS VDD clk n218 n183 n883 n217 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_3_ VSS VDD clk n216 n183 n980 n215 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_2_ VSS VDD clk n214 n183 n946 n213 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_1_ VSS VDD clk n212 n183 n941 n211 ASYNC_DFFHx1_ASAP7_75t_R
Xsum2_reg_0_ VSS VDD clk n210 n183 n868 n209 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_12_ VSS VDD clk n208 n183 n919 n207 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_11_ VSS VDD clk n206 n183 n900 n205 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_10_ VSS VDD clk n204 n183 n943 n203 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_9_ VSS VDD clk n202 n183 n882 n201 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_8_ VSS VDD clk n200 n183 n928 n199 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_7_ VSS VDD clk n198 n183 n926 n197 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_6_ VSS VDD clk n196 n183 n886 n195 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_5_ VSS VDD clk n194 n183 n888 n193 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_4_ VSS VDD clk n192 n183 n937 n191 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_3_ VSS VDD clk n190 n183 n929 n189 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_2_ VSS VDD clk n188 n183 n1009 n187 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_1_ VSS VDD clk n186 n183 n907 n185 ASYNC_DFFHx1_ASAP7_75t_R
Xsum3_reg_0_ VSS VDD clk n184 n183 n901 n182 ASYNC_DFFHx1_ASAP7_75t_R
XU940 VSS VDD n345 n1057 BUFx10_ASAP7_75t_R
XU908 VSS VDD n253 n1046 BUFx3_ASAP7_75t_R
XU909 VSS VDD n279 n1045 BUFx3_ASAP7_75t_R
XU910 VSS VDD n201 n1048 BUFx3_ASAP7_75t_R
XU911 VSS VDD n227 n1047 BUFx3_ASAP7_75t_R
XU1139 VSS VDD n223 n1031 BUFx5_ASAP7_75t_R
XU1140 VSS VDD n263 n1027 BUFx5_ASAP7_75t_R
XU1141 VSS VDD n241 n1029 BUFx5_ASAP7_75t_R
XU1208 VSS VDD n197 n1035 BUFx5_ASAP7_75t_R
XU1210 VSS VDD n249 n1028 BUFx5_ASAP7_75t_R
XU1212 VSS VDD n275 n1025 BUFx5_ASAP7_75t_R
XU1214 VSS VDD n237 n1030 BUFx5_ASAP7_75t_R
XU1216 VSS VDD n211 n1034 BUFx5_ASAP7_75t_R
XU1218 VSS VDD n185 n1037 BUFx5_ASAP7_75t_R
XU1220 VSS VDD n215 n1033 BUFx5_ASAP7_75t_R
XU1222 VSS VDD n219 n1032 BUFx5_ASAP7_75t_R
XU1224 VSS VDD n189 n1036 BUFx5_ASAP7_75t_R
XU1226 VSS VDD n267 n1026 BUFx5_ASAP7_75t_R
XU1230 VSS VDD n193 n1276 BUFx5_ASAP7_75t_R
XU1232 VSS VDD n245 n1258 BUFx5_ASAP7_75t_R
XU1234 VSS VDD n271 n1249 BUFx5_ASAP7_75t_R
Xin_data1_dff_reg_127_ VSS VDD clk n857 in_data1_dff[127] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_126_ VSS VDD clk n856 in_data1_dff[126] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_125_ VSS VDD clk n855 in_data1_dff[125] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_124_ VSS VDD clk n854 in_data1_dff[124] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_123_ VSS VDD clk n853 in_data1_dff[123] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_122_ VSS VDD clk n852 in_data1_dff[122] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_121_ VSS VDD clk n851 in_data1_dff[121] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_120_ VSS VDD clk n850 in_data1_dff[120] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_119_ VSS VDD clk n849 in_data1_dff[119] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_118_ VSS VDD clk n848 in_data1_dff[118] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_117_ VSS VDD clk n847 in_data1_dff[117] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_116_ VSS VDD clk n846 in_data1_dff[116] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_115_ VSS VDD clk n845 in_data1_dff[115] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_114_ VSS VDD clk n844 in_data1_dff[114] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_113_ VSS VDD clk n843 in_data1_dff[113] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_112_ VSS VDD clk n842 in_data1_dff[112] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_111_ VSS VDD clk n841 in_data1_dff[111] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_110_ VSS VDD clk n840 in_data1_dff[110] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_109_ VSS VDD clk n839 in_data1_dff[109] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_108_ VSS VDD clk n838 in_data1_dff[108] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_107_ VSS VDD clk n837 in_data1_dff[107] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_106_ VSS VDD clk n836 in_data1_dff[106] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_105_ VSS VDD clk n835 in_data1_dff[105] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_104_ VSS VDD clk n834 in_data1_dff[104] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_103_ VSS VDD clk n833 in_data1_dff[103] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_102_ VSS VDD clk n832 in_data1_dff[102] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_101_ VSS VDD clk n831 in_data1_dff[101] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_100_ VSS VDD clk n830 in_data1_dff[100] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_99_ VSS VDD clk n829 in_data1_dff[99] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_98_ VSS VDD clk n828 in_data1_dff[98] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_97_ VSS VDD clk n827 in_data1_dff[97] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_96_ VSS VDD clk n826 in_data1_dff[96] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_95_ VSS VDD clk n825 in_data1_dff[95] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_94_ VSS VDD clk n824 in_data1_dff[94] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_93_ VSS VDD clk n823 in_data1_dff[93] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_92_ VSS VDD clk n822 in_data1_dff[92] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_91_ VSS VDD clk n821 in_data1_dff[91] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_90_ VSS VDD clk n820 in_data1_dff[90] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_89_ VSS VDD clk n819 in_data1_dff[89] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_88_ VSS VDD clk n818 in_data1_dff[88] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_87_ VSS VDD clk n817 in_data1_dff[87] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_86_ VSS VDD clk n816 in_data1_dff[86] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_85_ VSS VDD clk n815 in_data1_dff[85] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_84_ VSS VDD clk n814 in_data1_dff[84] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_83_ VSS VDD clk n813 in_data1_dff[83] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_82_ VSS VDD clk n812 in_data1_dff[82] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_81_ VSS VDD clk n811 in_data1_dff[81] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_80_ VSS VDD clk n810 in_data1_dff[80] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_79_ VSS VDD clk n809 in_data1_dff[79] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_78_ VSS VDD clk n808 in_data1_dff[78] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_77_ VSS VDD clk n807 in_data1_dff[77] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_76_ VSS VDD clk n806 in_data1_dff[76] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_75_ VSS VDD clk n805 in_data1_dff[75] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_74_ VSS VDD clk n804 in_data1_dff[74] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_73_ VSS VDD clk n803 in_data1_dff[73] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_72_ VSS VDD clk n802 in_data1_dff[72] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_71_ VSS VDD clk n801 in_data1_dff[71] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_70_ VSS VDD clk n800 in_data1_dff[70] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_69_ VSS VDD clk n799 in_data1_dff[69] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_68_ VSS VDD clk n798 in_data1_dff[68] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_67_ VSS VDD clk n797 in_data1_dff[67] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_66_ VSS VDD clk n796 in_data1_dff[66] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_65_ VSS VDD clk n795 in_data1_dff[65] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_64_ VSS VDD clk n794 in_data1_dff[64] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_63_ VSS VDD clk n793 in_data1_dff[63] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_62_ VSS VDD clk n792 in_data1_dff[62] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_61_ VSS VDD clk n791 in_data1_dff[61] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_60_ VSS VDD clk n790 in_data1_dff[60] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_59_ VSS VDD clk n789 in_data1_dff[59] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_58_ VSS VDD clk n788 in_data1_dff[58] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_57_ VSS VDD clk n787 in_data1_dff[57] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_56_ VSS VDD clk n786 in_data1_dff[56] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_55_ VSS VDD clk n785 in_data1_dff[55] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_54_ VSS VDD clk n784 in_data1_dff[54] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_53_ VSS VDD clk n783 in_data1_dff[53] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_52_ VSS VDD clk n782 in_data1_dff[52] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_51_ VSS VDD clk n781 in_data1_dff[51] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_50_ VSS VDD clk n780 in_data1_dff[50] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_49_ VSS VDD clk n779 in_data1_dff[49] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_48_ VSS VDD clk n778 in_data1_dff[48] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_47_ VSS VDD clk n777 in_data1_dff[47] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_46_ VSS VDD clk n776 in_data1_dff[46] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_45_ VSS VDD clk n775 in_data1_dff[45] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_44_ VSS VDD clk n774 in_data1_dff[44] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_43_ VSS VDD clk n773 in_data1_dff[43] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_42_ VSS VDD clk n772 in_data1_dff[42] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_41_ VSS VDD clk n771 in_data1_dff[41] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_40_ VSS VDD clk n770 in_data1_dff[40] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_39_ VSS VDD clk n769 in_data1_dff[39] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_38_ VSS VDD clk n768 in_data1_dff[38] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_37_ VSS VDD clk n767 in_data1_dff[37] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_36_ VSS VDD clk n766 in_data1_dff[36] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_35_ VSS VDD clk n765 in_data1_dff[35] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_34_ VSS VDD clk n764 in_data1_dff[34] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_33_ VSS VDD clk n763 in_data1_dff[33] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_32_ VSS VDD clk n762 in_data1_dff[32] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_31_ VSS VDD clk n761 in_data1_dff[31] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_30_ VSS VDD clk n760 in_data1_dff[30] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_29_ VSS VDD clk n759 in_data1_dff[29] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_28_ VSS VDD clk n758 in_data1_dff[28] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_27_ VSS VDD clk n757 in_data1_dff[27] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_26_ VSS VDD clk n756 in_data1_dff[26] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_25_ VSS VDD clk n755 in_data1_dff[25] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_24_ VSS VDD clk n754 in_data1_dff[24] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_23_ VSS VDD clk n753 in_data1_dff[23] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_22_ VSS VDD clk n752 in_data1_dff[22] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_21_ VSS VDD clk n751 in_data1_dff[21] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_20_ VSS VDD clk n750 in_data1_dff[20] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_19_ VSS VDD clk n749 in_data1_dff[19] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_18_ VSS VDD clk n748 in_data1_dff[18] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_17_ VSS VDD clk n747 in_data1_dff[17] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_16_ VSS VDD clk n746 in_data1_dff[16] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_15_ VSS VDD clk n745 in_data1_dff[15] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_14_ VSS VDD clk n744 in_data1_dff[14] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_13_ VSS VDD clk n743 in_data1_dff[13] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_12_ VSS VDD clk n742 in_data1_dff[12] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_11_ VSS VDD clk n741 in_data1_dff[11] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_10_ VSS VDD clk n740 in_data1_dff[10] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_9_ VSS VDD clk n739 in_data1_dff[9] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_8_ VSS VDD clk n738 in_data1_dff[8] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_7_ VSS VDD clk n737 in_data1_dff[7] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_6_ VSS VDD clk n736 in_data1_dff[6] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_5_ VSS VDD clk n735 in_data1_dff[5] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_4_ VSS VDD clk n734 in_data1_dff[4] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_3_ VSS VDD clk n733 in_data1_dff[3] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_2_ VSS VDD clk n732 in_data1_dff[2] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_1_ VSS VDD clk n731 in_data1_dff[1] DFFHQNx1_ASAP7_75t_R
Xin_data1_dff_reg_0_ VSS VDD clk n730 in_data1_dff[0] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_127_ VSS VDD clk n729 in_data2_dff[127] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_126_ VSS VDD clk n728 in_data2_dff[126] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_125_ VSS VDD clk n727 in_data2_dff[125] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_124_ VSS VDD clk n726 in_data2_dff[124] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_123_ VSS VDD clk n725 in_data2_dff[123] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_122_ VSS VDD clk n724 in_data2_dff[122] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_121_ VSS VDD clk n723 in_data2_dff[121] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_120_ VSS VDD clk n722 in_data2_dff[120] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_119_ VSS VDD clk n721 in_data2_dff[119] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_118_ VSS VDD clk n720 in_data2_dff[118] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_117_ VSS VDD clk n719 in_data2_dff[117] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_116_ VSS VDD clk n718 in_data2_dff[116] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_115_ VSS VDD clk n717 in_data2_dff[115] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_114_ VSS VDD clk n716 in_data2_dff[114] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_113_ VSS VDD clk n715 in_data2_dff[113] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_112_ VSS VDD clk n714 in_data2_dff[112] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_111_ VSS VDD clk n713 in_data2_dff[111] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_110_ VSS VDD clk n712 in_data2_dff[110] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_109_ VSS VDD clk n711 in_data2_dff[109] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_108_ VSS VDD clk n710 in_data2_dff[108] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_107_ VSS VDD clk n709 in_data2_dff[107] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_106_ VSS VDD clk n708 in_data2_dff[106] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_105_ VSS VDD clk n707 in_data2_dff[105] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_104_ VSS VDD clk n706 in_data2_dff[104] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_103_ VSS VDD clk n705 in_data2_dff[103] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_102_ VSS VDD clk n704 in_data2_dff[102] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_101_ VSS VDD clk n703 in_data2_dff[101] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_100_ VSS VDD clk n702 in_data2_dff[100] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_99_ VSS VDD clk n701 in_data2_dff[99] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_98_ VSS VDD clk n700 in_data2_dff[98] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_97_ VSS VDD clk n699 in_data2_dff[97] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_96_ VSS VDD clk n698 in_data2_dff[96] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_95_ VSS VDD clk n697 in_data2_dff[95] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_94_ VSS VDD clk n696 in_data2_dff[94] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_93_ VSS VDD clk n695 in_data2_dff[93] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_92_ VSS VDD clk n694 in_data2_dff[92] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_91_ VSS VDD clk n693 in_data2_dff[91] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_90_ VSS VDD clk n692 in_data2_dff[90] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_89_ VSS VDD clk n691 in_data2_dff[89] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_88_ VSS VDD clk n690 in_data2_dff[88] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_87_ VSS VDD clk n689 in_data2_dff[87] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_86_ VSS VDD clk n688 in_data2_dff[86] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_85_ VSS VDD clk n687 in_data2_dff[85] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_84_ VSS VDD clk n686 in_data2_dff[84] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_83_ VSS VDD clk n685 in_data2_dff[83] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_82_ VSS VDD clk n684 in_data2_dff[82] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_81_ VSS VDD clk n683 in_data2_dff[81] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_80_ VSS VDD clk n682 in_data2_dff[80] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_79_ VSS VDD clk n681 in_data2_dff[79] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_78_ VSS VDD clk n680 in_data2_dff[78] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_77_ VSS VDD clk n679 in_data2_dff[77] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_76_ VSS VDD clk n678 in_data2_dff[76] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_75_ VSS VDD clk n677 in_data2_dff[75] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_74_ VSS VDD clk n676 in_data2_dff[74] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_73_ VSS VDD clk n675 in_data2_dff[73] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_72_ VSS VDD clk n674 in_data2_dff[72] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_71_ VSS VDD clk n673 in_data2_dff[71] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_70_ VSS VDD clk n672 in_data2_dff[70] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_69_ VSS VDD clk n671 in_data2_dff[69] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_68_ VSS VDD clk n670 in_data2_dff[68] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_67_ VSS VDD clk n669 in_data2_dff[67] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_66_ VSS VDD clk n668 in_data2_dff[66] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_65_ VSS VDD clk n667 in_data2_dff[65] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_64_ VSS VDD clk n666 in_data2_dff[64] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_63_ VSS VDD clk n665 in_data2_dff[63] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_62_ VSS VDD clk n664 in_data2_dff[62] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_61_ VSS VDD clk n663 in_data2_dff[61] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_60_ VSS VDD clk n662 in_data2_dff[60] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_59_ VSS VDD clk n661 in_data2_dff[59] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_58_ VSS VDD clk n660 in_data2_dff[58] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_57_ VSS VDD clk n659 in_data2_dff[57] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_56_ VSS VDD clk n658 in_data2_dff[56] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_55_ VSS VDD clk n657 in_data2_dff[55] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_54_ VSS VDD clk n656 in_data2_dff[54] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_53_ VSS VDD clk n655 in_data2_dff[53] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_52_ VSS VDD clk n654 in_data2_dff[52] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_51_ VSS VDD clk n653 in_data2_dff[51] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_50_ VSS VDD clk n652 in_data2_dff[50] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_49_ VSS VDD clk n651 in_data2_dff[49] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_48_ VSS VDD clk n650 in_data2_dff[48] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_47_ VSS VDD clk n649 in_data2_dff[47] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_46_ VSS VDD clk n648 in_data2_dff[46] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_45_ VSS VDD clk n647 in_data2_dff[45] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_44_ VSS VDD clk n646 in_data2_dff[44] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_43_ VSS VDD clk n645 in_data2_dff[43] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_42_ VSS VDD clk n644 in_data2_dff[42] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_41_ VSS VDD clk n643 in_data2_dff[41] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_40_ VSS VDD clk n642 in_data2_dff[40] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_39_ VSS VDD clk n641 in_data2_dff[39] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_38_ VSS VDD clk n640 in_data2_dff[38] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_37_ VSS VDD clk n639 in_data2_dff[37] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_36_ VSS VDD clk n638 in_data2_dff[36] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_35_ VSS VDD clk n637 in_data2_dff[35] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_34_ VSS VDD clk n636 in_data2_dff[34] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_33_ VSS VDD clk n635 in_data2_dff[33] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_32_ VSS VDD clk n634 in_data2_dff[32] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_31_ VSS VDD clk n633 in_data2_dff[31] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_30_ VSS VDD clk n632 in_data2_dff[30] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_29_ VSS VDD clk n631 in_data2_dff[29] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_28_ VSS VDD clk n630 in_data2_dff[28] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_27_ VSS VDD clk n629 in_data2_dff[27] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_26_ VSS VDD clk n628 in_data2_dff[26] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_25_ VSS VDD clk n627 in_data2_dff[25] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_24_ VSS VDD clk n626 in_data2_dff[24] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_23_ VSS VDD clk n625 in_data2_dff[23] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_22_ VSS VDD clk n624 in_data2_dff[22] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_21_ VSS VDD clk n623 in_data2_dff[21] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_20_ VSS VDD clk n622 in_data2_dff[20] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_19_ VSS VDD clk n621 in_data2_dff[19] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_18_ VSS VDD clk n620 in_data2_dff[18] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_17_ VSS VDD clk n619 in_data2_dff[17] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_16_ VSS VDD clk n618 in_data2_dff[16] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_15_ VSS VDD clk n617 in_data2_dff[15] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_14_ VSS VDD clk n616 in_data2_dff[14] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_13_ VSS VDD clk n615 in_data2_dff[13] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_12_ VSS VDD clk n614 in_data2_dff[12] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_11_ VSS VDD clk n613 in_data2_dff[11] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_10_ VSS VDD clk n612 in_data2_dff[10] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_9_ VSS VDD clk n611 in_data2_dff[9] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_8_ VSS VDD clk n610 in_data2_dff[8] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_7_ VSS VDD clk n609 in_data2_dff[7] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_6_ VSS VDD clk n608 in_data2_dff[6] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_5_ VSS VDD clk n607 in_data2_dff[5] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_4_ VSS VDD clk n606 in_data2_dff[4] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_3_ VSS VDD clk n605 in_data2_dff[3] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_2_ VSS VDD clk n604 in_data2_dff[2] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_1_ VSS VDD clk n603 in_data2_dff[1] DFFHQNx1_ASAP7_75t_R
Xin_data2_dff_reg_0_ VSS VDD clk n602 in_data2_dff[0] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_127_ VSS VDD clk n601 in_data3_dff[127] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_126_ VSS VDD clk n600 in_data3_dff[126] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_125_ VSS VDD clk n599 in_data3_dff[125] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_124_ VSS VDD clk n598 in_data3_dff[124] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_123_ VSS VDD clk n597 in_data3_dff[123] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_122_ VSS VDD clk n596 in_data3_dff[122] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_121_ VSS VDD clk n595 in_data3_dff[121] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_120_ VSS VDD clk n594 in_data3_dff[120] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_119_ VSS VDD clk n593 in_data3_dff[119] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_118_ VSS VDD clk n592 in_data3_dff[118] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_117_ VSS VDD clk n591 in_data3_dff[117] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_116_ VSS VDD clk n590 in_data3_dff[116] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_115_ VSS VDD clk n589 in_data3_dff[115] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_114_ VSS VDD clk n588 in_data3_dff[114] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_113_ VSS VDD clk n587 in_data3_dff[113] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_112_ VSS VDD clk n586 in_data3_dff[112] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_111_ VSS VDD clk n585 in_data3_dff[111] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_110_ VSS VDD clk n584 in_data3_dff[110] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_109_ VSS VDD clk n583 in_data3_dff[109] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_108_ VSS VDD clk n582 in_data3_dff[108] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_107_ VSS VDD clk n581 in_data3_dff[107] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_106_ VSS VDD clk n580 in_data3_dff[106] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_105_ VSS VDD clk n579 in_data3_dff[105] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_104_ VSS VDD clk n578 in_data3_dff[104] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_103_ VSS VDD clk n577 in_data3_dff[103] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_102_ VSS VDD clk n576 in_data3_dff[102] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_101_ VSS VDD clk n575 in_data3_dff[101] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_100_ VSS VDD clk n574 in_data3_dff[100] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_99_ VSS VDD clk n573 in_data3_dff[99] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_98_ VSS VDD clk n572 in_data3_dff[98] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_97_ VSS VDD clk n571 in_data3_dff[97] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_96_ VSS VDD clk n570 in_data3_dff[96] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_95_ VSS VDD clk n569 in_data3_dff[95] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_94_ VSS VDD clk n568 in_data3_dff[94] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_93_ VSS VDD clk n567 in_data3_dff[93] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_92_ VSS VDD clk n566 in_data3_dff[92] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_91_ VSS VDD clk n565 in_data3_dff[91] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_90_ VSS VDD clk n564 in_data3_dff[90] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_89_ VSS VDD clk n563 in_data3_dff[89] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_88_ VSS VDD clk n562 in_data3_dff[88] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_87_ VSS VDD clk n561 in_data3_dff[87] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_86_ VSS VDD clk n560 in_data3_dff[86] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_85_ VSS VDD clk n559 in_data3_dff[85] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_84_ VSS VDD clk n558 in_data3_dff[84] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_83_ VSS VDD clk n557 in_data3_dff[83] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_82_ VSS VDD clk n556 in_data3_dff[82] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_81_ VSS VDD clk n555 in_data3_dff[81] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_80_ VSS VDD clk n554 in_data3_dff[80] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_79_ VSS VDD clk n553 in_data3_dff[79] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_78_ VSS VDD clk n552 in_data3_dff[78] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_77_ VSS VDD clk n551 in_data3_dff[77] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_76_ VSS VDD clk n550 in_data3_dff[76] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_75_ VSS VDD clk n549 in_data3_dff[75] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_74_ VSS VDD clk n548 in_data3_dff[74] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_73_ VSS VDD clk n547 in_data3_dff[73] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_72_ VSS VDD clk n546 in_data3_dff[72] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_71_ VSS VDD clk n545 in_data3_dff[71] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_70_ VSS VDD clk n544 in_data3_dff[70] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_69_ VSS VDD clk n543 in_data3_dff[69] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_68_ VSS VDD clk n542 in_data3_dff[68] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_67_ VSS VDD clk n541 in_data3_dff[67] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_66_ VSS VDD clk n540 in_data3_dff[66] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_65_ VSS VDD clk n539 in_data3_dff[65] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_64_ VSS VDD clk n538 in_data3_dff[64] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_63_ VSS VDD clk n537 in_data3_dff[63] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_62_ VSS VDD clk n536 in_data3_dff[62] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_61_ VSS VDD clk n535 in_data3_dff[61] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_60_ VSS VDD clk n534 in_data3_dff[60] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_59_ VSS VDD clk n533 in_data3_dff[59] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_58_ VSS VDD clk n532 in_data3_dff[58] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_57_ VSS VDD clk n531 in_data3_dff[57] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_56_ VSS VDD clk n530 in_data3_dff[56] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_55_ VSS VDD clk n529 in_data3_dff[55] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_54_ VSS VDD clk n528 in_data3_dff[54] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_53_ VSS VDD clk n527 in_data3_dff[53] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_52_ VSS VDD clk n526 in_data3_dff[52] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_51_ VSS VDD clk n525 in_data3_dff[51] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_50_ VSS VDD clk n524 in_data3_dff[50] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_49_ VSS VDD clk n523 in_data3_dff[49] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_48_ VSS VDD clk n522 in_data3_dff[48] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_47_ VSS VDD clk n521 in_data3_dff[47] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_46_ VSS VDD clk n520 in_data3_dff[46] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_45_ VSS VDD clk n519 in_data3_dff[45] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_44_ VSS VDD clk n518 in_data3_dff[44] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_43_ VSS VDD clk n517 in_data3_dff[43] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_42_ VSS VDD clk n516 in_data3_dff[42] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_41_ VSS VDD clk n515 in_data3_dff[41] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_40_ VSS VDD clk n514 in_data3_dff[40] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_39_ VSS VDD clk n513 in_data3_dff[39] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_38_ VSS VDD clk n512 in_data3_dff[38] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_37_ VSS VDD clk n511 in_data3_dff[37] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_36_ VSS VDD clk n510 in_data3_dff[36] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_35_ VSS VDD clk n509 in_data3_dff[35] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_34_ VSS VDD clk n508 in_data3_dff[34] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_33_ VSS VDD clk n507 in_data3_dff[33] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_32_ VSS VDD clk n506 in_data3_dff[32] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_31_ VSS VDD clk n505 in_data3_dff[31] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_30_ VSS VDD clk n504 in_data3_dff[30] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_29_ VSS VDD clk n503 in_data3_dff[29] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_28_ VSS VDD clk n502 in_data3_dff[28] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_27_ VSS VDD clk n501 in_data3_dff[27] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_26_ VSS VDD clk n500 in_data3_dff[26] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_25_ VSS VDD clk n499 in_data3_dff[25] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_24_ VSS VDD clk n498 in_data3_dff[24] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_23_ VSS VDD clk n497 in_data3_dff[23] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_22_ VSS VDD clk n496 in_data3_dff[22] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_21_ VSS VDD clk n495 in_data3_dff[21] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_20_ VSS VDD clk n494 in_data3_dff[20] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_19_ VSS VDD clk n493 in_data3_dff[19] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_18_ VSS VDD clk n492 in_data3_dff[18] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_17_ VSS VDD clk n491 in_data3_dff[17] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_16_ VSS VDD clk n490 in_data3_dff[16] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_15_ VSS VDD clk n489 in_data3_dff[15] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_14_ VSS VDD clk n488 in_data3_dff[14] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_13_ VSS VDD clk n487 in_data3_dff[13] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_12_ VSS VDD clk n486 in_data3_dff[12] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_11_ VSS VDD clk n485 in_data3_dff[11] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_10_ VSS VDD clk n484 in_data3_dff[10] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_9_ VSS VDD clk n483 in_data3_dff[9] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_8_ VSS VDD clk n482 in_data3_dff[8] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_7_ VSS VDD clk n481 in_data3_dff[7] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_6_ VSS VDD clk n480 in_data3_dff[6] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_5_ VSS VDD clk n479 in_data3_dff[5] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_4_ VSS VDD clk n478 in_data3_dff[4] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_3_ VSS VDD clk n477 in_data3_dff[3] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_2_ VSS VDD clk n476 in_data3_dff[2] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_1_ VSS VDD clk n475 in_data3_dff[1] DFFHQNx1_ASAP7_75t_R
Xin_data3_dff_reg_0_ VSS VDD clk n474 in_data3_dff[0] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_127_ VSS VDD clk n473 in_data4_dff[127] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_126_ VSS VDD clk n472 in_data4_dff[126] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_125_ VSS VDD clk n471 in_data4_dff[125] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_124_ VSS VDD clk n470 in_data4_dff[124] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_123_ VSS VDD clk n469 in_data4_dff[123] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_122_ VSS VDD clk n468 in_data4_dff[122] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_121_ VSS VDD clk n467 in_data4_dff[121] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_120_ VSS VDD clk n466 in_data4_dff[120] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_119_ VSS VDD clk n465 in_data4_dff[119] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_118_ VSS VDD clk n464 in_data4_dff[118] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_117_ VSS VDD clk n463 in_data4_dff[117] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_116_ VSS VDD clk n462 in_data4_dff[116] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_115_ VSS VDD clk n461 in_data4_dff[115] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_114_ VSS VDD clk n460 in_data4_dff[114] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_113_ VSS VDD clk n459 in_data4_dff[113] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_112_ VSS VDD clk n458 in_data4_dff[112] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_111_ VSS VDD clk n457 in_data4_dff[111] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_110_ VSS VDD clk n456 in_data4_dff[110] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_109_ VSS VDD clk n455 in_data4_dff[109] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_108_ VSS VDD clk n454 in_data4_dff[108] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_107_ VSS VDD clk n453 in_data4_dff[107] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_106_ VSS VDD clk n452 in_data4_dff[106] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_105_ VSS VDD clk n451 in_data4_dff[105] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_104_ VSS VDD clk n450 in_data4_dff[104] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_103_ VSS VDD clk n449 in_data4_dff[103] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_102_ VSS VDD clk n448 in_data4_dff[102] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_101_ VSS VDD clk n447 in_data4_dff[101] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_100_ VSS VDD clk n446 in_data4_dff[100] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_99_ VSS VDD clk n445 in_data4_dff[99] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_98_ VSS VDD clk n444 in_data4_dff[98] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_97_ VSS VDD clk n443 in_data4_dff[97] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_96_ VSS VDD clk n442 in_data4_dff[96] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_95_ VSS VDD clk n441 in_data4_dff[95] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_94_ VSS VDD clk n440 in_data4_dff[94] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_93_ VSS VDD clk n439 in_data4_dff[93] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_92_ VSS VDD clk n438 in_data4_dff[92] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_91_ VSS VDD clk n437 in_data4_dff[91] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_90_ VSS VDD clk n436 in_data4_dff[90] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_89_ VSS VDD clk n435 in_data4_dff[89] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_88_ VSS VDD clk n434 in_data4_dff[88] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_87_ VSS VDD clk n433 in_data4_dff[87] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_86_ VSS VDD clk n432 in_data4_dff[86] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_85_ VSS VDD clk n431 in_data4_dff[85] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_84_ VSS VDD clk n430 in_data4_dff[84] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_83_ VSS VDD clk n429 in_data4_dff[83] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_82_ VSS VDD clk n428 in_data4_dff[82] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_81_ VSS VDD clk n427 in_data4_dff[81] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_80_ VSS VDD clk n426 in_data4_dff[80] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_79_ VSS VDD clk n425 in_data4_dff[79] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_78_ VSS VDD clk n424 in_data4_dff[78] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_77_ VSS VDD clk n423 in_data4_dff[77] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_76_ VSS VDD clk n422 in_data4_dff[76] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_75_ VSS VDD clk n421 in_data4_dff[75] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_74_ VSS VDD clk n420 in_data4_dff[74] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_73_ VSS VDD clk n419 in_data4_dff[73] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_72_ VSS VDD clk n418 in_data4_dff[72] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_71_ VSS VDD clk n417 in_data4_dff[71] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_70_ VSS VDD clk n416 in_data4_dff[70] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_69_ VSS VDD clk n415 in_data4_dff[69] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_68_ VSS VDD clk n414 in_data4_dff[68] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_67_ VSS VDD clk n413 in_data4_dff[67] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_66_ VSS VDD clk n412 in_data4_dff[66] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_65_ VSS VDD clk n411 in_data4_dff[65] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_64_ VSS VDD clk n410 in_data4_dff[64] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_63_ VSS VDD clk n409 in_data4_dff[63] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_62_ VSS VDD clk n408 in_data4_dff[62] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_61_ VSS VDD clk n407 in_data4_dff[61] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_60_ VSS VDD clk n406 in_data4_dff[60] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_59_ VSS VDD clk n405 in_data4_dff[59] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_58_ VSS VDD clk n404 in_data4_dff[58] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_57_ VSS VDD clk n403 in_data4_dff[57] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_56_ VSS VDD clk n402 in_data4_dff[56] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_55_ VSS VDD clk n401 in_data4_dff[55] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_54_ VSS VDD clk n400 in_data4_dff[54] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_53_ VSS VDD clk n399 in_data4_dff[53] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_52_ VSS VDD clk n398 in_data4_dff[52] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_51_ VSS VDD clk n397 in_data4_dff[51] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_50_ VSS VDD clk n396 in_data4_dff[50] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_49_ VSS VDD clk n395 in_data4_dff[49] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_48_ VSS VDD clk n394 in_data4_dff[48] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_47_ VSS VDD clk n393 in_data4_dff[47] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_46_ VSS VDD clk n392 in_data4_dff[46] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_45_ VSS VDD clk n391 in_data4_dff[45] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_44_ VSS VDD clk n390 in_data4_dff[44] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_43_ VSS VDD clk n389 in_data4_dff[43] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_42_ VSS VDD clk n388 in_data4_dff[42] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_41_ VSS VDD clk n387 in_data4_dff[41] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_40_ VSS VDD clk n386 in_data4_dff[40] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_39_ VSS VDD clk n385 in_data4_dff[39] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_38_ VSS VDD clk n384 in_data4_dff[38] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_37_ VSS VDD clk n383 in_data4_dff[37] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_36_ VSS VDD clk n382 in_data4_dff[36] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_35_ VSS VDD clk n381 in_data4_dff[35] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_34_ VSS VDD clk n380 in_data4_dff[34] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_33_ VSS VDD clk n379 in_data4_dff[33] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_32_ VSS VDD clk n378 in_data4_dff[32] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_31_ VSS VDD clk n377 in_data4_dff[31] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_30_ VSS VDD clk n376 in_data4_dff[30] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_29_ VSS VDD clk n375 in_data4_dff[29] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_28_ VSS VDD clk n374 in_data4_dff[28] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_27_ VSS VDD clk n373 in_data4_dff[27] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_26_ VSS VDD clk n372 in_data4_dff[26] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_25_ VSS VDD clk n371 in_data4_dff[25] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_24_ VSS VDD clk n370 in_data4_dff[24] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_23_ VSS VDD clk n369 in_data4_dff[23] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_22_ VSS VDD clk n368 in_data4_dff[22] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_21_ VSS VDD clk n367 in_data4_dff[21] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_20_ VSS VDD clk n366 in_data4_dff[20] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_19_ VSS VDD clk n365 in_data4_dff[19] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_18_ VSS VDD clk n364 in_data4_dff[18] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_17_ VSS VDD clk n363 in_data4_dff[17] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_16_ VSS VDD clk n362 in_data4_dff[16] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_15_ VSS VDD clk n361 in_data4_dff[15] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_14_ VSS VDD clk n360 in_data4_dff[14] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_13_ VSS VDD clk n359 in_data4_dff[13] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_12_ VSS VDD clk n358 in_data4_dff[12] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_11_ VSS VDD clk n357 in_data4_dff[11] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_10_ VSS VDD clk n356 in_data4_dff[10] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_9_ VSS VDD clk n355 in_data4_dff[9] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_8_ VSS VDD clk n354 in_data4_dff[8] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_7_ VSS VDD clk n353 in_data4_dff[7] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_6_ VSS VDD clk n352 in_data4_dff[6] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_5_ VSS VDD clk n351 in_data4_dff[5] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_4_ VSS VDD clk n350 in_data4_dff[4] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_3_ VSS VDD clk n349 in_data4_dff[3] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_2_ VSS VDD clk n348 in_data4_dff[2] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_1_ VSS VDD clk n347 in_data4_dff[1] DFFHQNx1_ASAP7_75t_R
Xin_data4_dff_reg_0_ VSS VDD clk n346 in_data4_dff[0] DFFHQNx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U243 VSS VDD in_data4_dff[120] in_data4_dff[96] in_data4_dff[88] DP_OP_657J1_125_1759_n332 DP_OP_657J1_125_1759_n333 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U242 VSS VDD in_data4_dff[80] in_data4_dff[72] in_data4_dff[64] DP_OP_657J1_125_1759_n330 DP_OP_657J1_125_1759_n331 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U241 VSS VDD in_data4_dff[56] in_data4_dff[48] in_data4_dff[40] DP_OP_657J1_125_1759_n328 DP_OP_657J1_125_1759_n329 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U240 VSS VDD in_data4_dff[32] in_data4_dff[24] in_data4_dff[16] DP_OP_657J1_125_1759_n326 DP_OP_657J1_125_1759_n327 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U239 VSS VDD in_data4_dff[8] in_data4_dff[0] in_data4_dff[4] DP_OP_657J1_125_1759_n324 DP_OP_657J1_125_1759_n325 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U238 VSS VDD in_data4_dff[12] in_data4_dff[20] in_data4_dff[28] DP_OP_657J1_125_1759_n322 DP_OP_657J1_125_1759_n323 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U237 VSS VDD in_data4_dff[36] in_data4_dff[44] in_data4_dff[52] DP_OP_657J1_125_1759_n320 DP_OP_657J1_125_1759_n321 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U236 VSS VDD in_data4_dff[60] in_data4_dff[68] in_data4_dff[76] DP_OP_657J1_125_1759_n318 DP_OP_657J1_125_1759_n319 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U235 VSS VDD in_data4_dff[84] in_data4_dff[124] in_data4_dff[92] DP_OP_657J1_125_1759_n316 DP_OP_657J1_125_1759_n317 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U234 VSS VDD in_data4_dff[100] in_data4_dff[116] in_data4_dff[108] DP_OP_657J1_125_1759_n314 DP_OP_657J1_125_1759_n315 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U232 VSS VDD DP_OP_657J1_125_1759_n317 DP_OP_657J1_125_1759_n311 DP_OP_657J1_125_1759_n319 DP_OP_657J1_125_1759_n312 DP_OP_657J1_125_1759_n313 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U231 VSS VDD DP_OP_657J1_125_1759_n315 DP_OP_657J1_125_1759_n321 DP_OP_657J1_125_1759_n323 DP_OP_657J1_125_1759_n309 DP_OP_657J1_125_1759_n310 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U230 VSS VDD DP_OP_657J1_125_1759_n325 DP_OP_657J1_125_1759_n327 DP_OP_657J1_125_1759_n329 DP_OP_657J1_125_1759_n307 DP_OP_657J1_125_1759_n308 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U228 VSS VDD DP_OP_657J1_125_1759_n331 DP_OP_657J1_125_1759_n333 DP_OP_657J1_125_1759_n304 DP_OP_657J1_125_1759_n305 DP_OP_657J1_125_1759_n306 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U225 VSS VDD in_data4_dff[105] in_data4_dff[97] in_data4_dff[89] DP_OP_657J1_125_1759_n300 DP_OP_657J1_125_1759_n301 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U224 VSS VDD in_data4_dff[81] in_data4_dff[73] in_data4_dff[65] DP_OP_657J1_125_1759_n298 DP_OP_657J1_125_1759_n299 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U223 VSS VDD in_data4_dff[57] in_data4_dff[49] in_data4_dff[41] DP_OP_657J1_125_1759_n296 DP_OP_657J1_125_1759_n297 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U222 VSS VDD in_data4_dff[33] in_data4_dff[25] in_data4_dff[17] DP_OP_657J1_125_1759_n294 DP_OP_657J1_125_1759_n295 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U221 VSS VDD in_data4_dff[9] in_data4_dff[45] in_data4_dff[125] DP_OP_657J1_125_1759_n292 DP_OP_657J1_125_1759_n293 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U220 VSS VDD in_data4_dff[1] in_data4_dff[37] in_data4_dff[5] DP_OP_657J1_125_1759_n290 DP_OP_657J1_125_1759_n291 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U219 VSS VDD in_data4_dff[117] in_data4_dff[61] in_data4_dff[109] DP_OP_657J1_125_1759_n288 DP_OP_657J1_125_1759_n289 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U218 VSS VDD in_data4_dff[13] in_data4_dff[29] in_data4_dff[101] DP_OP_657J1_125_1759_n286 DP_OP_657J1_125_1759_n287 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U217 VSS VDD in_data4_dff[21] in_data4_dff[93] in_data4_dff[53] DP_OP_657J1_125_1759_n284 DP_OP_657J1_125_1759_n285 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U216 VSS VDD in_data4_dff[69] in_data4_dff[85] in_data4_dff[77] DP_OP_657J1_125_1759_n282 DP_OP_657J1_125_1759_n283 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U214 VSS VDD DP_OP_657J1_125_1759_n332 DP_OP_657J1_125_1759_n279 DP_OP_657J1_125_1759_n330 DP_OP_657J1_125_1759_n280 DP_OP_657J1_125_1759_n281 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U212 VSS VDD DP_OP_657J1_125_1759_n328 DP_OP_657J1_125_1759_n316 DP_OP_657J1_125_1759_n276 DP_OP_657J1_125_1759_n277 DP_OP_657J1_125_1759_n278 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U211 VSS VDD DP_OP_657J1_125_1759_n318 DP_OP_657J1_125_1759_n314 DP_OP_657J1_125_1759_n320 DP_OP_657J1_125_1759_n274 DP_OP_657J1_125_1759_n275 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U210 VSS VDD DP_OP_657J1_125_1759_n322 DP_OP_657J1_125_1759_n324 DP_OP_657J1_125_1759_n326 DP_OP_657J1_125_1759_n272 DP_OP_657J1_125_1759_n273 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U209 VSS VDD DP_OP_657J1_125_1759_n293 DP_OP_657J1_125_1759_n283 DP_OP_657J1_125_1759_n295 DP_OP_657J1_125_1759_n270 DP_OP_657J1_125_1759_n271 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U208 VSS VDD DP_OP_657J1_125_1759_n291 DP_OP_657J1_125_1759_n285 DP_OP_657J1_125_1759_n289 DP_OP_657J1_125_1759_n268 DP_OP_657J1_125_1759_n269 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U207 VSS VDD DP_OP_657J1_125_1759_n299 DP_OP_657J1_125_1759_n287 DP_OP_657J1_125_1759_n297 DP_OP_657J1_125_1759_n266 DP_OP_657J1_125_1759_n267 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U205 VSS VDD DP_OP_657J1_125_1759_n312 DP_OP_657J1_125_1759_n281 DP_OP_657J1_125_1759_n263 DP_OP_657J1_125_1759_n264 DP_OP_657J1_125_1759_n265 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U204 VSS VDD DP_OP_657J1_125_1759_n273 DP_OP_657J1_125_1759_n275 DP_OP_657J1_125_1759_n278 DP_OP_657J1_125_1759_n261 DP_OP_657J1_125_1759_n262 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U203 VSS VDD DP_OP_657J1_125_1759_n307 DP_OP_657J1_125_1759_n309 DP_OP_657J1_125_1759_n271 DP_OP_657J1_125_1759_n259 DP_OP_657J1_125_1759_n260 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U201 VSS VDD DP_OP_657J1_125_1759_n267 DP_OP_657J1_125_1759_n269 DP_OP_657J1_125_1759_n256 DP_OP_657J1_125_1759_n257 DP_OP_657J1_125_1759_n258 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U199 VSS VDD DP_OP_657J1_125_1759_n260 DP_OP_657J1_125_1759_n262 DP_OP_657J1_125_1759_n253 DP_OP_657J1_125_1759_n254 DP_OP_657J1_125_1759_n255 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U195 VSS VDD in_data4_dff[106] in_data4_dff[98] in_data4_dff[90] DP_OP_657J1_125_1759_n248 DP_OP_657J1_125_1759_n249 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U194 VSS VDD in_data4_dff[82] in_data4_dff[74] in_data4_dff[66] DP_OP_657J1_125_1759_n246 DP_OP_657J1_125_1759_n247 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U193 VSS VDD in_data4_dff[126] in_data4_dff[22] in_data4_dff[118] DP_OP_657J1_125_1759_n244 DP_OP_657J1_125_1759_n245 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U192 VSS VDD in_data4_dff[58] in_data4_dff[110] in_data4_dff[50] DP_OP_657J1_125_1759_n242 DP_OP_657J1_125_1759_n243 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U191 VSS VDD in_data4_dff[42] in_data4_dff[102] in_data4_dff[94] DP_OP_657J1_125_1759_n240 DP_OP_657J1_125_1759_n241 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U190 VSS VDD in_data4_dff[34] in_data4_dff[6] in_data4_dff[26] DP_OP_657J1_125_1759_n238 DP_OP_657J1_125_1759_n239 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U189 VSS VDD in_data4_dff[18] in_data4_dff[86] in_data4_dff[10] DP_OP_657J1_125_1759_n236 DP_OP_657J1_125_1759_n237 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U188 VSS VDD in_data4_dff[2] in_data4_dff[78] in_data4_dff[14] DP_OP_657J1_125_1759_n234 DP_OP_657J1_125_1759_n235 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U187 VSS VDD in_data4_dff[70] in_data4_dff[38] in_data4_dff[62] DP_OP_657J1_125_1759_n232 DP_OP_657J1_125_1759_n233 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U186 VSS VDD in_data4_dff[30] in_data4_dff[54] in_data4_dff[46] DP_OP_657J1_125_1759_n230 DP_OP_657J1_125_1759_n231 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U184 VSS VDD DP_OP_657J1_125_1759_n300 DP_OP_657J1_125_1759_n227 DP_OP_657J1_125_1759_n298 DP_OP_657J1_125_1759_n228 DP_OP_657J1_125_1759_n229 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U182 VSS VDD DP_OP_657J1_125_1759_n296 DP_OP_657J1_125_1759_n282 DP_OP_657J1_125_1759_n224 DP_OP_657J1_125_1759_n225 DP_OP_657J1_125_1759_n226 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U181 VSS VDD DP_OP_657J1_125_1759_n294 DP_OP_657J1_125_1759_n290 DP_OP_657J1_125_1759_n284 DP_OP_657J1_125_1759_n222 DP_OP_657J1_125_1759_n223 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U180 VSS VDD DP_OP_657J1_125_1759_n292 DP_OP_657J1_125_1759_n286 DP_OP_657J1_125_1759_n288 DP_OP_657J1_125_1759_n220 DP_OP_657J1_125_1759_n221 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U178 VSS VDD DP_OP_657J1_125_1759_n274 DP_OP_657J1_125_1759_n280 DP_OP_657J1_125_1759_n217 DP_OP_657J1_125_1759_n218 DP_OP_657J1_125_1759_n219 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U176 VSS VDD DP_OP_657J1_125_1759_n243 DP_OP_657J1_125_1759_n235 DP_OP_657J1_125_1759_n214 DP_OP_657J1_125_1759_n215 DP_OP_657J1_125_1759_n216 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U175 VSS VDD DP_OP_657J1_125_1759_n247 DP_OP_657J1_125_1759_n237 DP_OP_657J1_125_1759_n249 DP_OP_657J1_125_1759_n212 DP_OP_657J1_125_1759_n213 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U174 VSS VDD DP_OP_657J1_125_1759_n245 DP_OP_657J1_125_1759_n233 DP_OP_657J1_125_1759_n239 DP_OP_657J1_125_1759_n210 DP_OP_657J1_125_1759_n211 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U172 VSS VDD DP_OP_657J1_125_1759_n277 DP_OP_657J1_125_1759_n229 DP_OP_657J1_125_1759_n207 DP_OP_657J1_125_1759_n208 DP_OP_657J1_125_1759_n209 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U171 VSS VDD DP_OP_657J1_125_1759_n223 DP_OP_657J1_125_1759_n221 DP_OP_657J1_125_1759_n226 DP_OP_657J1_125_1759_n205 DP_OP_657J1_125_1759_n206 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U170 VSS VDD DP_OP_657J1_125_1759_n266 DP_OP_657J1_125_1759_n270 DP_OP_657J1_125_1759_n268 DP_OP_657J1_125_1759_n203 DP_OP_657J1_125_1759_n204 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U168 VSS VDD DP_OP_657J1_125_1759_n261 DP_OP_657J1_125_1759_n264 DP_OP_657J1_125_1759_n200 DP_OP_657J1_125_1759_n201 DP_OP_657J1_125_1759_n202 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U166 VSS VDD DP_OP_657J1_125_1759_n213 DP_OP_657J1_125_1759_n211 DP_OP_657J1_125_1759_n197 DP_OP_657J1_125_1759_n198 DP_OP_657J1_125_1759_n199 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U165 VSS VDD DP_OP_657J1_125_1759_n259 DP_OP_657J1_125_1759_n209 DP_OP_657J1_125_1759_n204 DP_OP_657J1_125_1759_n195 DP_OP_657J1_125_1759_n196 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U164 VSS VDD DP_OP_657J1_125_1759_n257 DP_OP_657J1_125_1759_n206 DP_OP_657J1_125_1759_n199 DP_OP_657J1_125_1759_n193 DP_OP_657J1_125_1759_n194 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U163 VSS VDD DP_OP_657J1_125_1759_n254 DP_OP_657J1_125_1759_n202 DP_OP_657J1_125_1759_n196 DP_OP_657J1_125_1759_n191 DP_OP_657J1_125_1759_n192 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U159 VSS VDD in_data4_dff[107] in_data4_dff[99] in_data4_dff[91] DP_OP_657J1_125_1759_n186 DP_OP_657J1_125_1759_n187 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U158 VSS VDD in_data4_dff[83] in_data4_dff[15] in_data4_dff[75] DP_OP_657J1_125_1759_n184 DP_OP_657J1_125_1759_n185 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U157 VSS VDD in_data4_dff[67] in_data4_dff[127] in_data4_dff[59] DP_OP_657J1_125_1759_n182 DP_OP_657J1_125_1759_n183 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U156 VSS VDD in_data4_dff[51] in_data4_dff[31] in_data4_dff[119] DP_OP_657J1_125_1759_n180 DP_OP_657J1_125_1759_n181 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U155 VSS VDD in_data4_dff[111] in_data4_dff[23] in_data4_dff[43] DP_OP_657J1_125_1759_n178 DP_OP_657J1_125_1759_n179 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U154 VSS VDD in_data4_dff[35] in_data4_dff[103] in_data4_dff[27] DP_OP_657J1_125_1759_n176 DP_OP_657J1_125_1759_n177 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U153 VSS VDD in_data4_dff[19] in_data4_dff[95] in_data4_dff[11] DP_OP_657J1_125_1759_n174 DP_OP_657J1_125_1759_n175 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U152 VSS VDD in_data4_dff[3] in_data4_dff[87] in_data4_dff[7] DP_OP_657J1_125_1759_n172 DP_OP_657J1_125_1759_n173 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U151 VSS VDD in_data4_dff[39] in_data4_dff[79] in_data4_dff[47] DP_OP_657J1_125_1759_n170 DP_OP_657J1_125_1759_n171 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U150 VSS VDD in_data4_dff[55] in_data4_dff[71] in_data4_dff[63] DP_OP_657J1_125_1759_n168 DP_OP_657J1_125_1759_n169 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U148 VSS VDD DP_OP_657J1_125_1759_n248 DP_OP_657J1_125_1759_n165 DP_OP_657J1_125_1759_n246 DP_OP_657J1_125_1759_n166 DP_OP_657J1_125_1759_n167 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U146 VSS VDD DP_OP_657J1_125_1759_n244 DP_OP_657J1_125_1759_n230 DP_OP_657J1_125_1759_n162 DP_OP_657J1_125_1759_n163 DP_OP_657J1_125_1759_n164 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U145 VSS VDD DP_OP_657J1_125_1759_n242 DP_OP_657J1_125_1759_n238 DP_OP_657J1_125_1759_n232 DP_OP_657J1_125_1759_n160 DP_OP_657J1_125_1759_n161 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U144 VSS VDD DP_OP_657J1_125_1759_n240 DP_OP_657J1_125_1759_n236 DP_OP_657J1_125_1759_n234 DP_OP_657J1_125_1759_n158 DP_OP_657J1_125_1759_n159 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U142 VSS VDD DP_OP_657J1_125_1759_n222 DP_OP_657J1_125_1759_n228 DP_OP_657J1_125_1759_n155 DP_OP_657J1_125_1759_n156 DP_OP_657J1_125_1759_n157 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U140 VSS VDD DP_OP_657J1_125_1759_n183 DP_OP_657J1_125_1759_n169 DP_OP_657J1_125_1759_n152 DP_OP_657J1_125_1759_n153 DP_OP_657J1_125_1759_n154 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U139 VSS VDD DP_OP_657J1_125_1759_n181 DP_OP_657J1_125_1759_n175 DP_OP_657J1_125_1759_n179 DP_OP_657J1_125_1759_n150 DP_OP_657J1_125_1759_n151 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U138 VSS VDD DP_OP_657J1_125_1759_n185 DP_OP_657J1_125_1759_n187 DP_OP_657J1_125_1759_n177 DP_OP_657J1_125_1759_n148 DP_OP_657J1_125_1759_n149 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U136 VSS VDD DP_OP_657J1_125_1759_n225 DP_OP_657J1_125_1759_n167 DP_OP_657J1_125_1759_n145 DP_OP_657J1_125_1759_n146 DP_OP_657J1_125_1759_n147 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U134 VSS VDD DP_OP_657J1_125_1759_n215 DP_OP_657J1_125_1759_n212 DP_OP_657J1_125_1759_n142 DP_OP_657J1_125_1759_n143 DP_OP_657J1_125_1759_n144 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U133 VSS VDD DP_OP_657J1_125_1759_n161 DP_OP_657J1_125_1759_n210 DP_OP_657J1_125_1759_n164 DP_OP_657J1_125_1759_n140 DP_OP_657J1_125_1759_n141 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U131 VSS VDD DP_OP_657J1_125_1759_n149 DP_OP_657J1_125_1759_n159 DP_OP_657J1_125_1759_n137 DP_OP_657J1_125_1759_n138 DP_OP_657J1_125_1759_n139 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U129 VSS VDD DP_OP_657J1_125_1759_n203 DP_OP_657J1_125_1759_n157 DP_OP_657J1_125_1759_n134 DP_OP_657J1_125_1759_n135 DP_OP_657J1_125_1759_n136 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U127 VSS VDD DP_OP_657J1_125_1759_n205 DP_OP_657J1_125_1759_n147 DP_OP_657J1_125_1759_n131 DP_OP_657J1_125_1759_n132 DP_OP_657J1_125_1759_n133 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U125 VSS VDD DP_OP_657J1_125_1759_n144 DP_OP_657J1_125_1759_n141 DP_OP_657J1_125_1759_n128 DP_OP_657J1_125_1759_n129 DP_OP_657J1_125_1759_n130 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U123 VSS VDD DP_OP_657J1_125_1759_n139 DP_OP_657J1_125_1759_n198 DP_OP_657J1_125_1759_n125 DP_OP_657J1_125_1759_n126 DP_OP_657J1_125_1759_n127 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U122 VSS VDD DP_OP_657J1_125_1759_n133 DP_OP_657J1_125_1759_n136 DP_OP_657J1_125_1759_n193 DP_OP_657J1_125_1759_n123 DP_OP_657J1_125_1759_n124 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U120 VSS VDD DP_OP_657J1_125_1759_n127 DP_OP_657J1_125_1759_n130 DP_OP_657J1_125_1759_n120 DP_OP_657J1_125_1759_n121 DP_OP_657J1_125_1759_n122 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U114 VSS VDD DP_OP_657J1_125_1759_n184 DP_OP_657J1_125_1759_n170 DP_OP_657J1_125_1759_n182 DP_OP_657J1_125_1759_n113 DP_OP_657J1_125_1759_n114 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U113 VSS VDD DP_OP_657J1_125_1759_n180 DP_OP_657J1_125_1759_n176 DP_OP_657J1_125_1759_n168 DP_OP_657J1_125_1759_n111 DP_OP_657J1_125_1759_n112 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U112 VSS VDD DP_OP_657J1_125_1759_n172 DP_OP_657J1_125_1759_n174 DP_OP_657J1_125_1759_n178 DP_OP_657J1_125_1759_n109 DP_OP_657J1_125_1759_n110 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U111 VSS VDD DP_OP_657J1_125_1759_n158 DP_OP_657J1_125_1759_n166 DP_OP_657J1_125_1759_n163 DP_OP_657J1_125_1759_n107 DP_OP_657J1_125_1759_n108 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U110 VSS VDD DP_OP_657J1_125_1759_n117 DP_OP_657J1_125_1759_n160 DP_OP_657J1_125_1759_n148 DP_OP_657J1_125_1759_n105 DP_OP_657J1_125_1759_n106 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U108 VSS VDD DP_OP_657J1_125_1759_n153 DP_OP_657J1_125_1759_n110 DP_OP_657J1_125_1759_n102 DP_OP_657J1_125_1759_n103 DP_OP_657J1_125_1759_n104 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U107 VSS VDD DP_OP_657J1_125_1759_n114 DP_OP_657J1_125_1759_n150 DP_OP_657J1_125_1759_n112 DP_OP_657J1_125_1759_n100 DP_OP_657J1_125_1759_n101 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U106 VSS VDD DP_OP_657J1_125_1759_n108 DP_OP_657J1_125_1759_n146 DP_OP_657J1_125_1759_n140 DP_OP_657J1_125_1759_n98 DP_OP_657J1_125_1759_n99 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U105 VSS VDD DP_OP_657J1_125_1759_n106 DP_OP_657J1_125_1759_n143 DP_OP_657J1_125_1759_n138 DP_OP_657J1_125_1759_n96 DP_OP_657J1_125_1759_n97 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U103 VSS VDD DP_OP_657J1_125_1759_n104 DP_OP_657J1_125_1759_n101 DP_OP_657J1_125_1759_n93 DP_OP_657J1_125_1759_n94 DP_OP_657J1_125_1759_n95 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U102 VSS VDD DP_OP_657J1_125_1759_n99 DP_OP_657J1_125_1759_n132 DP_OP_657J1_125_1759_n129 DP_OP_657J1_125_1759_n91 DP_OP_657J1_125_1759_n92 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U101 VSS VDD DP_OP_657J1_125_1759_n126 DP_OP_657J1_125_1759_n97 DP_OP_657J1_125_1759_n95 DP_OP_657J1_125_1759_n89 DP_OP_657J1_125_1759_n90 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U100 VSS VDD DP_OP_657J1_125_1759_n92 DP_OP_657J1_125_1759_n123 DP_OP_657J1_125_1759_n121 DP_OP_657J1_125_1759_n87 DP_OP_657J1_125_1759_n88 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U98 VSS VDD DP_OP_657J1_125_1759_n109 DP_OP_657J1_125_1759_n116 DP_OP_657J1_125_1759_n113 DP_OP_657J1_125_1759_n84 DP_OP_657J1_125_1759_n85 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U96 VSS VDD DP_OP_657J1_125_1759_n107 DP_OP_657J1_125_1759_n105 DP_OP_657J1_125_1759_n81 DP_OP_657J1_125_1759_n82 DP_OP_657J1_125_1759_n83 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U95 VSS VDD DP_OP_657J1_125_1759_n100 DP_OP_657J1_125_1759_n85 DP_OP_657J1_125_1759_n103 DP_OP_657J1_125_1759_n79 DP_OP_657J1_125_1759_n80 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U94 VSS VDD DP_OP_657J1_125_1759_n83 DP_OP_657J1_125_1759_n98 DP_OP_657J1_125_1759_n96 DP_OP_657J1_125_1759_n77 DP_OP_657J1_125_1759_n78 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U92 VSS VDD DP_OP_657J1_125_1759_n94 DP_OP_657J1_125_1759_n80 DP_OP_657J1_125_1759_n74 DP_OP_657J1_125_1759_n75 DP_OP_657J1_125_1759_n76 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U91 VSS VDD DP_OP_657J1_125_1759_n89 DP_OP_657J1_125_1759_n78 DP_OP_657J1_125_1759_n76 DP_OP_657J1_125_1759_n72 DP_OP_657J1_125_1759_n73 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U89 VSS VDD DP_OP_657J1_125_1759_n82 DP_OP_657J1_125_1759_n79 DP_OP_657J1_125_1759_n69 DP_OP_657J1_125_1759_n70 DP_OP_657J1_125_1759_n71 FAx1_ASAP7_75t_R
XDP_OP_657J1_125_1759_U88 VSS VDD DP_OP_657J1_125_1759_n71 DP_OP_657J1_125_1759_n77 DP_OP_657J1_125_1759_n75 DP_OP_657J1_125_1759_n67 DP_OP_657J1_125_1759_n68 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U243 VSS VDD in_data3_dff[120] in_data3_dff[96] in_data3_dff[88] DP_OP_656J1_124_1759_n332 DP_OP_656J1_124_1759_n333 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U242 VSS VDD in_data3_dff[80] in_data3_dff[72] in_data3_dff[64] DP_OP_656J1_124_1759_n330 DP_OP_656J1_124_1759_n331 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U241 VSS VDD in_data3_dff[56] in_data3_dff[48] in_data3_dff[40] DP_OP_656J1_124_1759_n328 DP_OP_656J1_124_1759_n329 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U240 VSS VDD in_data3_dff[32] in_data3_dff[24] in_data3_dff[16] DP_OP_656J1_124_1759_n326 DP_OP_656J1_124_1759_n327 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U239 VSS VDD in_data3_dff[8] in_data3_dff[0] in_data3_dff[4] DP_OP_656J1_124_1759_n324 DP_OP_656J1_124_1759_n325 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U238 VSS VDD in_data3_dff[12] in_data3_dff[20] in_data3_dff[28] DP_OP_656J1_124_1759_n322 DP_OP_656J1_124_1759_n323 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U237 VSS VDD in_data3_dff[36] in_data3_dff[44] in_data3_dff[52] DP_OP_656J1_124_1759_n320 DP_OP_656J1_124_1759_n321 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U236 VSS VDD in_data3_dff[60] in_data3_dff[68] in_data3_dff[76] DP_OP_656J1_124_1759_n318 DP_OP_656J1_124_1759_n319 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U235 VSS VDD in_data3_dff[84] in_data3_dff[124] in_data3_dff[92] DP_OP_656J1_124_1759_n316 DP_OP_656J1_124_1759_n317 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U234 VSS VDD in_data3_dff[100] in_data3_dff[116] in_data3_dff[108] DP_OP_656J1_124_1759_n314 DP_OP_656J1_124_1759_n315 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U232 VSS VDD DP_OP_656J1_124_1759_n317 DP_OP_656J1_124_1759_n311 DP_OP_656J1_124_1759_n319 DP_OP_656J1_124_1759_n312 DP_OP_656J1_124_1759_n313 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U231 VSS VDD DP_OP_656J1_124_1759_n315 DP_OP_656J1_124_1759_n321 DP_OP_656J1_124_1759_n323 DP_OP_656J1_124_1759_n309 DP_OP_656J1_124_1759_n310 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U230 VSS VDD DP_OP_656J1_124_1759_n325 DP_OP_656J1_124_1759_n327 DP_OP_656J1_124_1759_n329 DP_OP_656J1_124_1759_n307 DP_OP_656J1_124_1759_n308 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U228 VSS VDD DP_OP_656J1_124_1759_n331 DP_OP_656J1_124_1759_n333 DP_OP_656J1_124_1759_n304 DP_OP_656J1_124_1759_n305 DP_OP_656J1_124_1759_n306 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U225 VSS VDD in_data3_dff[105] in_data3_dff[97] in_data3_dff[89] DP_OP_656J1_124_1759_n300 DP_OP_656J1_124_1759_n301 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U224 VSS VDD in_data3_dff[81] in_data3_dff[73] in_data3_dff[65] DP_OP_656J1_124_1759_n298 DP_OP_656J1_124_1759_n299 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U223 VSS VDD in_data3_dff[57] in_data3_dff[49] in_data3_dff[41] DP_OP_656J1_124_1759_n296 DP_OP_656J1_124_1759_n297 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U222 VSS VDD in_data3_dff[33] in_data3_dff[25] in_data3_dff[17] DP_OP_656J1_124_1759_n294 DP_OP_656J1_124_1759_n295 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U221 VSS VDD in_data3_dff[9] in_data3_dff[45] in_data3_dff[125] DP_OP_656J1_124_1759_n292 DP_OP_656J1_124_1759_n293 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U220 VSS VDD in_data3_dff[1] in_data3_dff[37] in_data3_dff[5] DP_OP_656J1_124_1759_n290 DP_OP_656J1_124_1759_n291 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U219 VSS VDD in_data3_dff[117] in_data3_dff[61] in_data3_dff[109] DP_OP_656J1_124_1759_n288 DP_OP_656J1_124_1759_n289 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U218 VSS VDD in_data3_dff[13] in_data3_dff[29] in_data3_dff[101] DP_OP_656J1_124_1759_n286 DP_OP_656J1_124_1759_n287 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U217 VSS VDD in_data3_dff[21] in_data3_dff[93] in_data3_dff[53] DP_OP_656J1_124_1759_n284 DP_OP_656J1_124_1759_n285 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U216 VSS VDD in_data3_dff[69] in_data3_dff[85] in_data3_dff[77] DP_OP_656J1_124_1759_n282 DP_OP_656J1_124_1759_n283 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U214 VSS VDD DP_OP_656J1_124_1759_n332 DP_OP_656J1_124_1759_n279 DP_OP_656J1_124_1759_n330 DP_OP_656J1_124_1759_n280 DP_OP_656J1_124_1759_n281 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U212 VSS VDD DP_OP_656J1_124_1759_n328 DP_OP_656J1_124_1759_n316 DP_OP_656J1_124_1759_n276 DP_OP_656J1_124_1759_n277 DP_OP_656J1_124_1759_n278 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U211 VSS VDD DP_OP_656J1_124_1759_n318 DP_OP_656J1_124_1759_n314 DP_OP_656J1_124_1759_n320 DP_OP_656J1_124_1759_n274 DP_OP_656J1_124_1759_n275 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U210 VSS VDD DP_OP_656J1_124_1759_n322 DP_OP_656J1_124_1759_n324 DP_OP_656J1_124_1759_n326 DP_OP_656J1_124_1759_n272 DP_OP_656J1_124_1759_n273 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U209 VSS VDD DP_OP_656J1_124_1759_n293 DP_OP_656J1_124_1759_n283 DP_OP_656J1_124_1759_n295 DP_OP_656J1_124_1759_n270 DP_OP_656J1_124_1759_n271 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U208 VSS VDD DP_OP_656J1_124_1759_n291 DP_OP_656J1_124_1759_n285 DP_OP_656J1_124_1759_n289 DP_OP_656J1_124_1759_n268 DP_OP_656J1_124_1759_n269 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U207 VSS VDD DP_OP_656J1_124_1759_n299 DP_OP_656J1_124_1759_n287 DP_OP_656J1_124_1759_n297 DP_OP_656J1_124_1759_n266 DP_OP_656J1_124_1759_n267 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U205 VSS VDD DP_OP_656J1_124_1759_n312 DP_OP_656J1_124_1759_n281 DP_OP_656J1_124_1759_n263 DP_OP_656J1_124_1759_n264 DP_OP_656J1_124_1759_n265 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U204 VSS VDD DP_OP_656J1_124_1759_n273 DP_OP_656J1_124_1759_n275 DP_OP_656J1_124_1759_n278 DP_OP_656J1_124_1759_n261 DP_OP_656J1_124_1759_n262 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U203 VSS VDD DP_OP_656J1_124_1759_n307 DP_OP_656J1_124_1759_n309 DP_OP_656J1_124_1759_n271 DP_OP_656J1_124_1759_n259 DP_OP_656J1_124_1759_n260 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U201 VSS VDD DP_OP_656J1_124_1759_n267 DP_OP_656J1_124_1759_n269 DP_OP_656J1_124_1759_n256 DP_OP_656J1_124_1759_n257 DP_OP_656J1_124_1759_n258 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U199 VSS VDD DP_OP_656J1_124_1759_n260 DP_OP_656J1_124_1759_n262 DP_OP_656J1_124_1759_n253 DP_OP_656J1_124_1759_n254 DP_OP_656J1_124_1759_n255 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U195 VSS VDD in_data3_dff[106] in_data3_dff[98] in_data3_dff[90] DP_OP_656J1_124_1759_n248 DP_OP_656J1_124_1759_n249 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U194 VSS VDD in_data3_dff[82] in_data3_dff[74] in_data3_dff[66] DP_OP_656J1_124_1759_n246 DP_OP_656J1_124_1759_n247 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U193 VSS VDD in_data3_dff[126] in_data3_dff[22] in_data3_dff[118] DP_OP_656J1_124_1759_n244 DP_OP_656J1_124_1759_n245 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U192 VSS VDD in_data3_dff[58] in_data3_dff[110] in_data3_dff[50] DP_OP_656J1_124_1759_n242 DP_OP_656J1_124_1759_n243 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U191 VSS VDD in_data3_dff[42] in_data3_dff[102] in_data3_dff[94] DP_OP_656J1_124_1759_n240 DP_OP_656J1_124_1759_n241 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U190 VSS VDD in_data3_dff[34] in_data3_dff[6] in_data3_dff[26] DP_OP_656J1_124_1759_n238 DP_OP_656J1_124_1759_n239 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U189 VSS VDD in_data3_dff[18] in_data3_dff[86] in_data3_dff[10] DP_OP_656J1_124_1759_n236 DP_OP_656J1_124_1759_n237 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U188 VSS VDD in_data3_dff[2] in_data3_dff[78] in_data3_dff[14] DP_OP_656J1_124_1759_n234 DP_OP_656J1_124_1759_n235 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U187 VSS VDD in_data3_dff[70] in_data3_dff[38] in_data3_dff[62] DP_OP_656J1_124_1759_n232 DP_OP_656J1_124_1759_n233 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U186 VSS VDD in_data3_dff[30] in_data3_dff[54] in_data3_dff[46] DP_OP_656J1_124_1759_n230 DP_OP_656J1_124_1759_n231 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U184 VSS VDD DP_OP_656J1_124_1759_n300 DP_OP_656J1_124_1759_n227 DP_OP_656J1_124_1759_n298 DP_OP_656J1_124_1759_n228 DP_OP_656J1_124_1759_n229 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U182 VSS VDD DP_OP_656J1_124_1759_n296 DP_OP_656J1_124_1759_n282 DP_OP_656J1_124_1759_n224 DP_OP_656J1_124_1759_n225 DP_OP_656J1_124_1759_n226 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U181 VSS VDD DP_OP_656J1_124_1759_n294 DP_OP_656J1_124_1759_n290 DP_OP_656J1_124_1759_n284 DP_OP_656J1_124_1759_n222 DP_OP_656J1_124_1759_n223 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U180 VSS VDD DP_OP_656J1_124_1759_n292 DP_OP_656J1_124_1759_n286 DP_OP_656J1_124_1759_n288 DP_OP_656J1_124_1759_n220 DP_OP_656J1_124_1759_n221 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U178 VSS VDD DP_OP_656J1_124_1759_n274 DP_OP_656J1_124_1759_n280 DP_OP_656J1_124_1759_n217 DP_OP_656J1_124_1759_n218 DP_OP_656J1_124_1759_n219 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U176 VSS VDD DP_OP_656J1_124_1759_n243 DP_OP_656J1_124_1759_n235 DP_OP_656J1_124_1759_n214 DP_OP_656J1_124_1759_n215 DP_OP_656J1_124_1759_n216 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U175 VSS VDD DP_OP_656J1_124_1759_n247 DP_OP_656J1_124_1759_n237 DP_OP_656J1_124_1759_n249 DP_OP_656J1_124_1759_n212 DP_OP_656J1_124_1759_n213 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U174 VSS VDD DP_OP_656J1_124_1759_n245 DP_OP_656J1_124_1759_n233 DP_OP_656J1_124_1759_n239 DP_OP_656J1_124_1759_n210 DP_OP_656J1_124_1759_n211 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U172 VSS VDD DP_OP_656J1_124_1759_n277 DP_OP_656J1_124_1759_n229 DP_OP_656J1_124_1759_n207 DP_OP_656J1_124_1759_n208 DP_OP_656J1_124_1759_n209 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U171 VSS VDD DP_OP_656J1_124_1759_n223 DP_OP_656J1_124_1759_n221 DP_OP_656J1_124_1759_n226 DP_OP_656J1_124_1759_n205 DP_OP_656J1_124_1759_n206 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U170 VSS VDD DP_OP_656J1_124_1759_n266 DP_OP_656J1_124_1759_n270 DP_OP_656J1_124_1759_n268 DP_OP_656J1_124_1759_n203 DP_OP_656J1_124_1759_n204 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U168 VSS VDD DP_OP_656J1_124_1759_n261 DP_OP_656J1_124_1759_n264 DP_OP_656J1_124_1759_n200 DP_OP_656J1_124_1759_n201 DP_OP_656J1_124_1759_n202 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U166 VSS VDD DP_OP_656J1_124_1759_n213 DP_OP_656J1_124_1759_n211 DP_OP_656J1_124_1759_n197 DP_OP_656J1_124_1759_n198 DP_OP_656J1_124_1759_n199 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U165 VSS VDD DP_OP_656J1_124_1759_n259 DP_OP_656J1_124_1759_n209 DP_OP_656J1_124_1759_n204 DP_OP_656J1_124_1759_n195 DP_OP_656J1_124_1759_n196 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U164 VSS VDD DP_OP_656J1_124_1759_n257 DP_OP_656J1_124_1759_n206 DP_OP_656J1_124_1759_n199 DP_OP_656J1_124_1759_n193 DP_OP_656J1_124_1759_n194 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U163 VSS VDD DP_OP_656J1_124_1759_n254 DP_OP_656J1_124_1759_n202 DP_OP_656J1_124_1759_n196 DP_OP_656J1_124_1759_n191 DP_OP_656J1_124_1759_n192 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U159 VSS VDD in_data3_dff[107] in_data3_dff[99] in_data3_dff[91] DP_OP_656J1_124_1759_n186 DP_OP_656J1_124_1759_n187 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U158 VSS VDD in_data3_dff[83] in_data3_dff[15] in_data3_dff[75] DP_OP_656J1_124_1759_n184 DP_OP_656J1_124_1759_n185 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U157 VSS VDD in_data3_dff[67] in_data3_dff[127] in_data3_dff[59] DP_OP_656J1_124_1759_n182 DP_OP_656J1_124_1759_n183 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U156 VSS VDD in_data3_dff[51] in_data3_dff[31] in_data3_dff[119] DP_OP_656J1_124_1759_n180 DP_OP_656J1_124_1759_n181 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U155 VSS VDD in_data3_dff[111] in_data3_dff[23] in_data3_dff[43] DP_OP_656J1_124_1759_n178 DP_OP_656J1_124_1759_n179 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U154 VSS VDD in_data3_dff[35] in_data3_dff[103] in_data3_dff[27] DP_OP_656J1_124_1759_n176 DP_OP_656J1_124_1759_n177 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U153 VSS VDD in_data3_dff[19] in_data3_dff[95] in_data3_dff[11] DP_OP_656J1_124_1759_n174 DP_OP_656J1_124_1759_n175 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U152 VSS VDD in_data3_dff[3] in_data3_dff[87] in_data3_dff[7] DP_OP_656J1_124_1759_n172 DP_OP_656J1_124_1759_n173 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U151 VSS VDD in_data3_dff[39] in_data3_dff[79] in_data3_dff[47] DP_OP_656J1_124_1759_n170 DP_OP_656J1_124_1759_n171 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U150 VSS VDD in_data3_dff[55] in_data3_dff[71] in_data3_dff[63] DP_OP_656J1_124_1759_n168 DP_OP_656J1_124_1759_n169 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U148 VSS VDD DP_OP_656J1_124_1759_n248 DP_OP_656J1_124_1759_n165 DP_OP_656J1_124_1759_n246 DP_OP_656J1_124_1759_n166 DP_OP_656J1_124_1759_n167 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U146 VSS VDD DP_OP_656J1_124_1759_n244 DP_OP_656J1_124_1759_n230 DP_OP_656J1_124_1759_n162 DP_OP_656J1_124_1759_n163 DP_OP_656J1_124_1759_n164 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U145 VSS VDD DP_OP_656J1_124_1759_n242 DP_OP_656J1_124_1759_n238 DP_OP_656J1_124_1759_n232 DP_OP_656J1_124_1759_n160 DP_OP_656J1_124_1759_n161 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U144 VSS VDD DP_OP_656J1_124_1759_n240 DP_OP_656J1_124_1759_n236 DP_OP_656J1_124_1759_n234 DP_OP_656J1_124_1759_n158 DP_OP_656J1_124_1759_n159 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U142 VSS VDD DP_OP_656J1_124_1759_n222 DP_OP_656J1_124_1759_n228 DP_OP_656J1_124_1759_n155 DP_OP_656J1_124_1759_n156 DP_OP_656J1_124_1759_n157 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U140 VSS VDD DP_OP_656J1_124_1759_n183 DP_OP_656J1_124_1759_n169 DP_OP_656J1_124_1759_n152 DP_OP_656J1_124_1759_n153 DP_OP_656J1_124_1759_n154 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U139 VSS VDD DP_OP_656J1_124_1759_n181 DP_OP_656J1_124_1759_n175 DP_OP_656J1_124_1759_n179 DP_OP_656J1_124_1759_n150 DP_OP_656J1_124_1759_n151 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U138 VSS VDD DP_OP_656J1_124_1759_n185 DP_OP_656J1_124_1759_n187 DP_OP_656J1_124_1759_n177 DP_OP_656J1_124_1759_n148 DP_OP_656J1_124_1759_n149 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U136 VSS VDD DP_OP_656J1_124_1759_n225 DP_OP_656J1_124_1759_n167 DP_OP_656J1_124_1759_n145 DP_OP_656J1_124_1759_n146 DP_OP_656J1_124_1759_n147 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U134 VSS VDD DP_OP_656J1_124_1759_n215 DP_OP_656J1_124_1759_n212 DP_OP_656J1_124_1759_n142 DP_OP_656J1_124_1759_n143 DP_OP_656J1_124_1759_n144 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U133 VSS VDD DP_OP_656J1_124_1759_n161 DP_OP_656J1_124_1759_n210 DP_OP_656J1_124_1759_n164 DP_OP_656J1_124_1759_n140 DP_OP_656J1_124_1759_n141 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U131 VSS VDD DP_OP_656J1_124_1759_n149 DP_OP_656J1_124_1759_n159 DP_OP_656J1_124_1759_n137 DP_OP_656J1_124_1759_n138 DP_OP_656J1_124_1759_n139 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U129 VSS VDD DP_OP_656J1_124_1759_n203 DP_OP_656J1_124_1759_n157 DP_OP_656J1_124_1759_n134 DP_OP_656J1_124_1759_n135 DP_OP_656J1_124_1759_n136 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U127 VSS VDD DP_OP_656J1_124_1759_n205 DP_OP_656J1_124_1759_n147 DP_OP_656J1_124_1759_n131 DP_OP_656J1_124_1759_n132 DP_OP_656J1_124_1759_n133 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U125 VSS VDD DP_OP_656J1_124_1759_n144 DP_OP_656J1_124_1759_n141 DP_OP_656J1_124_1759_n128 DP_OP_656J1_124_1759_n129 DP_OP_656J1_124_1759_n130 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U123 VSS VDD DP_OP_656J1_124_1759_n139 DP_OP_656J1_124_1759_n198 DP_OP_656J1_124_1759_n125 DP_OP_656J1_124_1759_n126 DP_OP_656J1_124_1759_n127 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U122 VSS VDD DP_OP_656J1_124_1759_n133 DP_OP_656J1_124_1759_n136 DP_OP_656J1_124_1759_n193 DP_OP_656J1_124_1759_n123 DP_OP_656J1_124_1759_n124 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U120 VSS VDD DP_OP_656J1_124_1759_n127 DP_OP_656J1_124_1759_n130 DP_OP_656J1_124_1759_n120 DP_OP_656J1_124_1759_n121 DP_OP_656J1_124_1759_n122 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U114 VSS VDD DP_OP_656J1_124_1759_n184 DP_OP_656J1_124_1759_n170 DP_OP_656J1_124_1759_n182 DP_OP_656J1_124_1759_n113 DP_OP_656J1_124_1759_n114 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U113 VSS VDD DP_OP_656J1_124_1759_n180 DP_OP_656J1_124_1759_n176 DP_OP_656J1_124_1759_n168 DP_OP_656J1_124_1759_n111 DP_OP_656J1_124_1759_n112 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U112 VSS VDD DP_OP_656J1_124_1759_n172 DP_OP_656J1_124_1759_n174 DP_OP_656J1_124_1759_n178 DP_OP_656J1_124_1759_n109 DP_OP_656J1_124_1759_n110 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U111 VSS VDD DP_OP_656J1_124_1759_n158 DP_OP_656J1_124_1759_n166 DP_OP_656J1_124_1759_n163 DP_OP_656J1_124_1759_n107 DP_OP_656J1_124_1759_n108 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U110 VSS VDD DP_OP_656J1_124_1759_n117 DP_OP_656J1_124_1759_n160 DP_OP_656J1_124_1759_n148 DP_OP_656J1_124_1759_n105 DP_OP_656J1_124_1759_n106 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U108 VSS VDD DP_OP_656J1_124_1759_n153 DP_OP_656J1_124_1759_n110 DP_OP_656J1_124_1759_n102 DP_OP_656J1_124_1759_n103 DP_OP_656J1_124_1759_n104 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U107 VSS VDD DP_OP_656J1_124_1759_n114 DP_OP_656J1_124_1759_n150 DP_OP_656J1_124_1759_n112 DP_OP_656J1_124_1759_n100 DP_OP_656J1_124_1759_n101 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U106 VSS VDD DP_OP_656J1_124_1759_n108 DP_OP_656J1_124_1759_n146 DP_OP_656J1_124_1759_n140 DP_OP_656J1_124_1759_n98 DP_OP_656J1_124_1759_n99 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U105 VSS VDD DP_OP_656J1_124_1759_n106 DP_OP_656J1_124_1759_n143 DP_OP_656J1_124_1759_n138 DP_OP_656J1_124_1759_n96 DP_OP_656J1_124_1759_n97 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U103 VSS VDD DP_OP_656J1_124_1759_n104 DP_OP_656J1_124_1759_n101 DP_OP_656J1_124_1759_n93 DP_OP_656J1_124_1759_n94 DP_OP_656J1_124_1759_n95 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U102 VSS VDD DP_OP_656J1_124_1759_n99 DP_OP_656J1_124_1759_n132 DP_OP_656J1_124_1759_n129 DP_OP_656J1_124_1759_n91 DP_OP_656J1_124_1759_n92 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U101 VSS VDD DP_OP_656J1_124_1759_n126 DP_OP_656J1_124_1759_n97 DP_OP_656J1_124_1759_n95 DP_OP_656J1_124_1759_n89 DP_OP_656J1_124_1759_n90 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U100 VSS VDD DP_OP_656J1_124_1759_n92 DP_OP_656J1_124_1759_n123 DP_OP_656J1_124_1759_n121 DP_OP_656J1_124_1759_n87 DP_OP_656J1_124_1759_n88 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U98 VSS VDD DP_OP_656J1_124_1759_n109 DP_OP_656J1_124_1759_n116 DP_OP_656J1_124_1759_n113 DP_OP_656J1_124_1759_n84 DP_OP_656J1_124_1759_n85 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U96 VSS VDD DP_OP_656J1_124_1759_n107 DP_OP_656J1_124_1759_n105 DP_OP_656J1_124_1759_n81 DP_OP_656J1_124_1759_n82 DP_OP_656J1_124_1759_n83 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U95 VSS VDD DP_OP_656J1_124_1759_n100 DP_OP_656J1_124_1759_n85 DP_OP_656J1_124_1759_n103 DP_OP_656J1_124_1759_n79 DP_OP_656J1_124_1759_n80 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U94 VSS VDD DP_OP_656J1_124_1759_n83 DP_OP_656J1_124_1759_n98 DP_OP_656J1_124_1759_n96 DP_OP_656J1_124_1759_n77 DP_OP_656J1_124_1759_n78 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U92 VSS VDD DP_OP_656J1_124_1759_n94 DP_OP_656J1_124_1759_n80 DP_OP_656J1_124_1759_n74 DP_OP_656J1_124_1759_n75 DP_OP_656J1_124_1759_n76 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U91 VSS VDD DP_OP_656J1_124_1759_n89 DP_OP_656J1_124_1759_n78 DP_OP_656J1_124_1759_n76 DP_OP_656J1_124_1759_n72 DP_OP_656J1_124_1759_n73 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U89 VSS VDD DP_OP_656J1_124_1759_n82 DP_OP_656J1_124_1759_n79 DP_OP_656J1_124_1759_n69 DP_OP_656J1_124_1759_n70 DP_OP_656J1_124_1759_n71 FAx1_ASAP7_75t_R
XDP_OP_656J1_124_1759_U88 VSS VDD DP_OP_656J1_124_1759_n71 DP_OP_656J1_124_1759_n77 DP_OP_656J1_124_1759_n75 DP_OP_656J1_124_1759_n67 DP_OP_656J1_124_1759_n68 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U243 VSS VDD in_data2_dff[120] in_data2_dff[96] in_data2_dff[88] DP_OP_655J1_123_1759_n332 DP_OP_655J1_123_1759_n333 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U242 VSS VDD in_data2_dff[80] in_data2_dff[72] in_data2_dff[64] DP_OP_655J1_123_1759_n330 DP_OP_655J1_123_1759_n331 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U241 VSS VDD in_data2_dff[56] in_data2_dff[48] in_data2_dff[40] DP_OP_655J1_123_1759_n328 DP_OP_655J1_123_1759_n329 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U240 VSS VDD in_data2_dff[32] in_data2_dff[24] in_data2_dff[16] DP_OP_655J1_123_1759_n326 DP_OP_655J1_123_1759_n327 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U239 VSS VDD in_data2_dff[8] in_data2_dff[0] in_data2_dff[4] DP_OP_655J1_123_1759_n324 DP_OP_655J1_123_1759_n325 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U238 VSS VDD in_data2_dff[12] in_data2_dff[20] in_data2_dff[28] DP_OP_655J1_123_1759_n322 DP_OP_655J1_123_1759_n323 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U237 VSS VDD in_data2_dff[36] in_data2_dff[44] in_data2_dff[52] DP_OP_655J1_123_1759_n320 DP_OP_655J1_123_1759_n321 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U236 VSS VDD in_data2_dff[60] in_data2_dff[68] in_data2_dff[76] DP_OP_655J1_123_1759_n318 DP_OP_655J1_123_1759_n319 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U235 VSS VDD in_data2_dff[84] in_data2_dff[124] in_data2_dff[92] DP_OP_655J1_123_1759_n316 DP_OP_655J1_123_1759_n317 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U234 VSS VDD in_data2_dff[100] in_data2_dff[116] in_data2_dff[108] DP_OP_655J1_123_1759_n314 DP_OP_655J1_123_1759_n315 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U232 VSS VDD DP_OP_655J1_123_1759_n317 DP_OP_655J1_123_1759_n311 DP_OP_655J1_123_1759_n319 DP_OP_655J1_123_1759_n312 DP_OP_655J1_123_1759_n313 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U231 VSS VDD DP_OP_655J1_123_1759_n315 DP_OP_655J1_123_1759_n321 DP_OP_655J1_123_1759_n323 DP_OP_655J1_123_1759_n309 DP_OP_655J1_123_1759_n310 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U230 VSS VDD DP_OP_655J1_123_1759_n325 DP_OP_655J1_123_1759_n327 DP_OP_655J1_123_1759_n329 DP_OP_655J1_123_1759_n307 DP_OP_655J1_123_1759_n308 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U228 VSS VDD DP_OP_655J1_123_1759_n331 DP_OP_655J1_123_1759_n333 DP_OP_655J1_123_1759_n304 DP_OP_655J1_123_1759_n305 DP_OP_655J1_123_1759_n306 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U225 VSS VDD in_data2_dff[105] in_data2_dff[97] in_data2_dff[89] DP_OP_655J1_123_1759_n300 DP_OP_655J1_123_1759_n301 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U224 VSS VDD in_data2_dff[81] in_data2_dff[73] in_data2_dff[65] DP_OP_655J1_123_1759_n298 DP_OP_655J1_123_1759_n299 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U223 VSS VDD in_data2_dff[57] in_data2_dff[49] in_data2_dff[41] DP_OP_655J1_123_1759_n296 DP_OP_655J1_123_1759_n297 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U222 VSS VDD in_data2_dff[33] in_data2_dff[25] in_data2_dff[17] DP_OP_655J1_123_1759_n294 DP_OP_655J1_123_1759_n295 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U221 VSS VDD in_data2_dff[9] in_data2_dff[45] in_data2_dff[125] DP_OP_655J1_123_1759_n292 DP_OP_655J1_123_1759_n293 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U220 VSS VDD in_data2_dff[1] in_data2_dff[37] in_data2_dff[5] DP_OP_655J1_123_1759_n290 DP_OP_655J1_123_1759_n291 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U219 VSS VDD in_data2_dff[117] in_data2_dff[61] in_data2_dff[109] DP_OP_655J1_123_1759_n288 DP_OP_655J1_123_1759_n289 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U218 VSS VDD in_data2_dff[13] in_data2_dff[29] in_data2_dff[101] DP_OP_655J1_123_1759_n286 DP_OP_655J1_123_1759_n287 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U217 VSS VDD in_data2_dff[21] in_data2_dff[93] in_data2_dff[53] DP_OP_655J1_123_1759_n284 DP_OP_655J1_123_1759_n285 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U216 VSS VDD in_data2_dff[69] in_data2_dff[85] in_data2_dff[77] DP_OP_655J1_123_1759_n282 DP_OP_655J1_123_1759_n283 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U214 VSS VDD DP_OP_655J1_123_1759_n332 DP_OP_655J1_123_1759_n279 DP_OP_655J1_123_1759_n330 DP_OP_655J1_123_1759_n280 DP_OP_655J1_123_1759_n281 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U212 VSS VDD DP_OP_655J1_123_1759_n328 DP_OP_655J1_123_1759_n316 DP_OP_655J1_123_1759_n276 DP_OP_655J1_123_1759_n277 DP_OP_655J1_123_1759_n278 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U211 VSS VDD DP_OP_655J1_123_1759_n318 DP_OP_655J1_123_1759_n314 DP_OP_655J1_123_1759_n320 DP_OP_655J1_123_1759_n274 DP_OP_655J1_123_1759_n275 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U210 VSS VDD DP_OP_655J1_123_1759_n322 DP_OP_655J1_123_1759_n324 DP_OP_655J1_123_1759_n326 DP_OP_655J1_123_1759_n272 DP_OP_655J1_123_1759_n273 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U209 VSS VDD DP_OP_655J1_123_1759_n293 DP_OP_655J1_123_1759_n283 DP_OP_655J1_123_1759_n295 DP_OP_655J1_123_1759_n270 DP_OP_655J1_123_1759_n271 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U208 VSS VDD DP_OP_655J1_123_1759_n291 DP_OP_655J1_123_1759_n285 DP_OP_655J1_123_1759_n289 DP_OP_655J1_123_1759_n268 DP_OP_655J1_123_1759_n269 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U207 VSS VDD DP_OP_655J1_123_1759_n299 DP_OP_655J1_123_1759_n287 DP_OP_655J1_123_1759_n297 DP_OP_655J1_123_1759_n266 DP_OP_655J1_123_1759_n267 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U205 VSS VDD DP_OP_655J1_123_1759_n312 DP_OP_655J1_123_1759_n281 DP_OP_655J1_123_1759_n263 DP_OP_655J1_123_1759_n264 DP_OP_655J1_123_1759_n265 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U204 VSS VDD DP_OP_655J1_123_1759_n273 DP_OP_655J1_123_1759_n275 DP_OP_655J1_123_1759_n278 DP_OP_655J1_123_1759_n261 DP_OP_655J1_123_1759_n262 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U203 VSS VDD DP_OP_655J1_123_1759_n307 DP_OP_655J1_123_1759_n309 DP_OP_655J1_123_1759_n271 DP_OP_655J1_123_1759_n259 DP_OP_655J1_123_1759_n260 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U201 VSS VDD DP_OP_655J1_123_1759_n267 DP_OP_655J1_123_1759_n269 DP_OP_655J1_123_1759_n256 DP_OP_655J1_123_1759_n257 DP_OP_655J1_123_1759_n258 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U199 VSS VDD DP_OP_655J1_123_1759_n260 DP_OP_655J1_123_1759_n262 DP_OP_655J1_123_1759_n253 DP_OP_655J1_123_1759_n254 DP_OP_655J1_123_1759_n255 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U195 VSS VDD in_data2_dff[106] in_data2_dff[98] in_data2_dff[90] DP_OP_655J1_123_1759_n248 DP_OP_655J1_123_1759_n249 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U194 VSS VDD in_data2_dff[82] in_data2_dff[74] in_data2_dff[66] DP_OP_655J1_123_1759_n246 DP_OP_655J1_123_1759_n247 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U193 VSS VDD in_data2_dff[126] in_data2_dff[22] in_data2_dff[118] DP_OP_655J1_123_1759_n244 DP_OP_655J1_123_1759_n245 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U192 VSS VDD in_data2_dff[58] in_data2_dff[110] in_data2_dff[50] DP_OP_655J1_123_1759_n242 DP_OP_655J1_123_1759_n243 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U191 VSS VDD in_data2_dff[42] in_data2_dff[102] in_data2_dff[94] DP_OP_655J1_123_1759_n240 DP_OP_655J1_123_1759_n241 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U190 VSS VDD in_data2_dff[34] in_data2_dff[6] in_data2_dff[26] DP_OP_655J1_123_1759_n238 DP_OP_655J1_123_1759_n239 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U189 VSS VDD in_data2_dff[18] in_data2_dff[86] in_data2_dff[10] DP_OP_655J1_123_1759_n236 DP_OP_655J1_123_1759_n237 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U188 VSS VDD in_data2_dff[2] in_data2_dff[78] in_data2_dff[14] DP_OP_655J1_123_1759_n234 DP_OP_655J1_123_1759_n235 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U187 VSS VDD in_data2_dff[70] in_data2_dff[38] in_data2_dff[62] DP_OP_655J1_123_1759_n232 DP_OP_655J1_123_1759_n233 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U186 VSS VDD in_data2_dff[30] in_data2_dff[54] in_data2_dff[46] DP_OP_655J1_123_1759_n230 DP_OP_655J1_123_1759_n231 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U184 VSS VDD DP_OP_655J1_123_1759_n300 DP_OP_655J1_123_1759_n227 DP_OP_655J1_123_1759_n298 DP_OP_655J1_123_1759_n228 DP_OP_655J1_123_1759_n229 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U182 VSS VDD DP_OP_655J1_123_1759_n296 DP_OP_655J1_123_1759_n282 DP_OP_655J1_123_1759_n224 DP_OP_655J1_123_1759_n225 DP_OP_655J1_123_1759_n226 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U181 VSS VDD DP_OP_655J1_123_1759_n294 DP_OP_655J1_123_1759_n290 DP_OP_655J1_123_1759_n284 DP_OP_655J1_123_1759_n222 DP_OP_655J1_123_1759_n223 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U180 VSS VDD DP_OP_655J1_123_1759_n292 DP_OP_655J1_123_1759_n286 DP_OP_655J1_123_1759_n288 DP_OP_655J1_123_1759_n220 DP_OP_655J1_123_1759_n221 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U178 VSS VDD DP_OP_655J1_123_1759_n274 DP_OP_655J1_123_1759_n280 DP_OP_655J1_123_1759_n217 DP_OP_655J1_123_1759_n218 DP_OP_655J1_123_1759_n219 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U176 VSS VDD DP_OP_655J1_123_1759_n243 DP_OP_655J1_123_1759_n235 DP_OP_655J1_123_1759_n214 DP_OP_655J1_123_1759_n215 DP_OP_655J1_123_1759_n216 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U175 VSS VDD DP_OP_655J1_123_1759_n247 DP_OP_655J1_123_1759_n237 DP_OP_655J1_123_1759_n249 DP_OP_655J1_123_1759_n212 DP_OP_655J1_123_1759_n213 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U174 VSS VDD DP_OP_655J1_123_1759_n245 DP_OP_655J1_123_1759_n233 DP_OP_655J1_123_1759_n239 DP_OP_655J1_123_1759_n210 DP_OP_655J1_123_1759_n211 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U172 VSS VDD DP_OP_655J1_123_1759_n277 DP_OP_655J1_123_1759_n229 DP_OP_655J1_123_1759_n207 DP_OP_655J1_123_1759_n208 DP_OP_655J1_123_1759_n209 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U171 VSS VDD DP_OP_655J1_123_1759_n223 DP_OP_655J1_123_1759_n221 DP_OP_655J1_123_1759_n226 DP_OP_655J1_123_1759_n205 DP_OP_655J1_123_1759_n206 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U170 VSS VDD DP_OP_655J1_123_1759_n266 DP_OP_655J1_123_1759_n270 DP_OP_655J1_123_1759_n268 DP_OP_655J1_123_1759_n203 DP_OP_655J1_123_1759_n204 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U168 VSS VDD DP_OP_655J1_123_1759_n261 DP_OP_655J1_123_1759_n264 DP_OP_655J1_123_1759_n200 DP_OP_655J1_123_1759_n201 DP_OP_655J1_123_1759_n202 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U166 VSS VDD DP_OP_655J1_123_1759_n213 DP_OP_655J1_123_1759_n211 DP_OP_655J1_123_1759_n197 DP_OP_655J1_123_1759_n198 DP_OP_655J1_123_1759_n199 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U165 VSS VDD DP_OP_655J1_123_1759_n259 DP_OP_655J1_123_1759_n209 DP_OP_655J1_123_1759_n204 DP_OP_655J1_123_1759_n195 DP_OP_655J1_123_1759_n196 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U164 VSS VDD DP_OP_655J1_123_1759_n257 DP_OP_655J1_123_1759_n206 DP_OP_655J1_123_1759_n199 DP_OP_655J1_123_1759_n193 DP_OP_655J1_123_1759_n194 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U163 VSS VDD DP_OP_655J1_123_1759_n254 DP_OP_655J1_123_1759_n202 DP_OP_655J1_123_1759_n196 DP_OP_655J1_123_1759_n191 DP_OP_655J1_123_1759_n192 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U159 VSS VDD in_data2_dff[107] in_data2_dff[99] in_data2_dff[91] DP_OP_655J1_123_1759_n186 DP_OP_655J1_123_1759_n187 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U158 VSS VDD in_data2_dff[83] in_data2_dff[15] in_data2_dff[75] DP_OP_655J1_123_1759_n184 DP_OP_655J1_123_1759_n185 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U157 VSS VDD in_data2_dff[67] in_data2_dff[127] in_data2_dff[59] DP_OP_655J1_123_1759_n182 DP_OP_655J1_123_1759_n183 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U156 VSS VDD in_data2_dff[51] in_data2_dff[31] in_data2_dff[119] DP_OP_655J1_123_1759_n180 DP_OP_655J1_123_1759_n181 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U155 VSS VDD in_data2_dff[111] in_data2_dff[23] in_data2_dff[43] DP_OP_655J1_123_1759_n178 DP_OP_655J1_123_1759_n179 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U154 VSS VDD in_data2_dff[35] in_data2_dff[103] in_data2_dff[27] DP_OP_655J1_123_1759_n176 DP_OP_655J1_123_1759_n177 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U153 VSS VDD in_data2_dff[19] in_data2_dff[95] in_data2_dff[11] DP_OP_655J1_123_1759_n174 DP_OP_655J1_123_1759_n175 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U152 VSS VDD in_data2_dff[3] in_data2_dff[87] in_data2_dff[7] DP_OP_655J1_123_1759_n172 DP_OP_655J1_123_1759_n173 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U151 VSS VDD in_data2_dff[39] in_data2_dff[79] in_data2_dff[47] DP_OP_655J1_123_1759_n170 DP_OP_655J1_123_1759_n171 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U150 VSS VDD in_data2_dff[55] in_data2_dff[71] in_data2_dff[63] DP_OP_655J1_123_1759_n168 DP_OP_655J1_123_1759_n169 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U148 VSS VDD DP_OP_655J1_123_1759_n248 DP_OP_655J1_123_1759_n165 DP_OP_655J1_123_1759_n246 DP_OP_655J1_123_1759_n166 DP_OP_655J1_123_1759_n167 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U146 VSS VDD DP_OP_655J1_123_1759_n244 DP_OP_655J1_123_1759_n230 DP_OP_655J1_123_1759_n162 DP_OP_655J1_123_1759_n163 DP_OP_655J1_123_1759_n164 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U145 VSS VDD DP_OP_655J1_123_1759_n242 DP_OP_655J1_123_1759_n238 DP_OP_655J1_123_1759_n232 DP_OP_655J1_123_1759_n160 DP_OP_655J1_123_1759_n161 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U144 VSS VDD DP_OP_655J1_123_1759_n240 DP_OP_655J1_123_1759_n236 DP_OP_655J1_123_1759_n234 DP_OP_655J1_123_1759_n158 DP_OP_655J1_123_1759_n159 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U142 VSS VDD DP_OP_655J1_123_1759_n222 DP_OP_655J1_123_1759_n228 DP_OP_655J1_123_1759_n155 DP_OP_655J1_123_1759_n156 DP_OP_655J1_123_1759_n157 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U140 VSS VDD DP_OP_655J1_123_1759_n183 DP_OP_655J1_123_1759_n169 DP_OP_655J1_123_1759_n152 DP_OP_655J1_123_1759_n153 DP_OP_655J1_123_1759_n154 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U139 VSS VDD DP_OP_655J1_123_1759_n181 DP_OP_655J1_123_1759_n175 DP_OP_655J1_123_1759_n179 DP_OP_655J1_123_1759_n150 DP_OP_655J1_123_1759_n151 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U138 VSS VDD DP_OP_655J1_123_1759_n185 DP_OP_655J1_123_1759_n187 DP_OP_655J1_123_1759_n177 DP_OP_655J1_123_1759_n148 DP_OP_655J1_123_1759_n149 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U136 VSS VDD DP_OP_655J1_123_1759_n225 DP_OP_655J1_123_1759_n167 DP_OP_655J1_123_1759_n145 DP_OP_655J1_123_1759_n146 DP_OP_655J1_123_1759_n147 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U134 VSS VDD DP_OP_655J1_123_1759_n215 DP_OP_655J1_123_1759_n212 DP_OP_655J1_123_1759_n142 DP_OP_655J1_123_1759_n143 DP_OP_655J1_123_1759_n144 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U133 VSS VDD DP_OP_655J1_123_1759_n161 DP_OP_655J1_123_1759_n210 DP_OP_655J1_123_1759_n164 DP_OP_655J1_123_1759_n140 DP_OP_655J1_123_1759_n141 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U131 VSS VDD DP_OP_655J1_123_1759_n149 DP_OP_655J1_123_1759_n159 DP_OP_655J1_123_1759_n137 DP_OP_655J1_123_1759_n138 DP_OP_655J1_123_1759_n139 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U129 VSS VDD DP_OP_655J1_123_1759_n203 DP_OP_655J1_123_1759_n157 DP_OP_655J1_123_1759_n134 DP_OP_655J1_123_1759_n135 DP_OP_655J1_123_1759_n136 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U127 VSS VDD DP_OP_655J1_123_1759_n205 DP_OP_655J1_123_1759_n147 DP_OP_655J1_123_1759_n131 DP_OP_655J1_123_1759_n132 DP_OP_655J1_123_1759_n133 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U125 VSS VDD DP_OP_655J1_123_1759_n144 DP_OP_655J1_123_1759_n141 DP_OP_655J1_123_1759_n128 DP_OP_655J1_123_1759_n129 DP_OP_655J1_123_1759_n130 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U123 VSS VDD DP_OP_655J1_123_1759_n139 DP_OP_655J1_123_1759_n198 DP_OP_655J1_123_1759_n125 DP_OP_655J1_123_1759_n126 DP_OP_655J1_123_1759_n127 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U122 VSS VDD DP_OP_655J1_123_1759_n133 DP_OP_655J1_123_1759_n136 DP_OP_655J1_123_1759_n193 DP_OP_655J1_123_1759_n123 DP_OP_655J1_123_1759_n124 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U120 VSS VDD DP_OP_655J1_123_1759_n127 DP_OP_655J1_123_1759_n130 DP_OP_655J1_123_1759_n120 DP_OP_655J1_123_1759_n121 DP_OP_655J1_123_1759_n122 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U114 VSS VDD DP_OP_655J1_123_1759_n184 DP_OP_655J1_123_1759_n170 DP_OP_655J1_123_1759_n182 DP_OP_655J1_123_1759_n113 DP_OP_655J1_123_1759_n114 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U113 VSS VDD DP_OP_655J1_123_1759_n180 DP_OP_655J1_123_1759_n176 DP_OP_655J1_123_1759_n168 DP_OP_655J1_123_1759_n111 DP_OP_655J1_123_1759_n112 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U112 VSS VDD DP_OP_655J1_123_1759_n172 DP_OP_655J1_123_1759_n174 DP_OP_655J1_123_1759_n178 DP_OP_655J1_123_1759_n109 DP_OP_655J1_123_1759_n110 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U111 VSS VDD DP_OP_655J1_123_1759_n158 DP_OP_655J1_123_1759_n166 DP_OP_655J1_123_1759_n163 DP_OP_655J1_123_1759_n107 DP_OP_655J1_123_1759_n108 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U110 VSS VDD DP_OP_655J1_123_1759_n117 DP_OP_655J1_123_1759_n160 DP_OP_655J1_123_1759_n148 DP_OP_655J1_123_1759_n105 DP_OP_655J1_123_1759_n106 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U108 VSS VDD DP_OP_655J1_123_1759_n153 DP_OP_655J1_123_1759_n110 DP_OP_655J1_123_1759_n102 DP_OP_655J1_123_1759_n103 DP_OP_655J1_123_1759_n104 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U107 VSS VDD DP_OP_655J1_123_1759_n114 DP_OP_655J1_123_1759_n150 DP_OP_655J1_123_1759_n112 DP_OP_655J1_123_1759_n100 DP_OP_655J1_123_1759_n101 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U106 VSS VDD DP_OP_655J1_123_1759_n108 DP_OP_655J1_123_1759_n146 DP_OP_655J1_123_1759_n140 DP_OP_655J1_123_1759_n98 DP_OP_655J1_123_1759_n99 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U105 VSS VDD DP_OP_655J1_123_1759_n106 DP_OP_655J1_123_1759_n143 DP_OP_655J1_123_1759_n138 DP_OP_655J1_123_1759_n96 DP_OP_655J1_123_1759_n97 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U103 VSS VDD DP_OP_655J1_123_1759_n104 DP_OP_655J1_123_1759_n101 DP_OP_655J1_123_1759_n93 DP_OP_655J1_123_1759_n94 DP_OP_655J1_123_1759_n95 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U102 VSS VDD DP_OP_655J1_123_1759_n99 DP_OP_655J1_123_1759_n132 DP_OP_655J1_123_1759_n129 DP_OP_655J1_123_1759_n91 DP_OP_655J1_123_1759_n92 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U101 VSS VDD DP_OP_655J1_123_1759_n126 DP_OP_655J1_123_1759_n97 DP_OP_655J1_123_1759_n95 DP_OP_655J1_123_1759_n89 DP_OP_655J1_123_1759_n90 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U100 VSS VDD DP_OP_655J1_123_1759_n92 DP_OP_655J1_123_1759_n123 DP_OP_655J1_123_1759_n121 DP_OP_655J1_123_1759_n87 DP_OP_655J1_123_1759_n88 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U98 VSS VDD DP_OP_655J1_123_1759_n109 DP_OP_655J1_123_1759_n116 DP_OP_655J1_123_1759_n113 DP_OP_655J1_123_1759_n84 DP_OP_655J1_123_1759_n85 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U96 VSS VDD DP_OP_655J1_123_1759_n107 DP_OP_655J1_123_1759_n105 DP_OP_655J1_123_1759_n81 DP_OP_655J1_123_1759_n82 DP_OP_655J1_123_1759_n83 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U95 VSS VDD DP_OP_655J1_123_1759_n100 DP_OP_655J1_123_1759_n85 DP_OP_655J1_123_1759_n103 DP_OP_655J1_123_1759_n79 DP_OP_655J1_123_1759_n80 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U94 VSS VDD DP_OP_655J1_123_1759_n83 DP_OP_655J1_123_1759_n98 DP_OP_655J1_123_1759_n96 DP_OP_655J1_123_1759_n77 DP_OP_655J1_123_1759_n78 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U92 VSS VDD DP_OP_655J1_123_1759_n94 DP_OP_655J1_123_1759_n80 DP_OP_655J1_123_1759_n74 DP_OP_655J1_123_1759_n75 DP_OP_655J1_123_1759_n76 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U91 VSS VDD DP_OP_655J1_123_1759_n89 DP_OP_655J1_123_1759_n78 DP_OP_655J1_123_1759_n76 DP_OP_655J1_123_1759_n72 DP_OP_655J1_123_1759_n73 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U89 VSS VDD DP_OP_655J1_123_1759_n82 DP_OP_655J1_123_1759_n79 DP_OP_655J1_123_1759_n69 DP_OP_655J1_123_1759_n70 DP_OP_655J1_123_1759_n71 FAx1_ASAP7_75t_R
XDP_OP_655J1_123_1759_U88 VSS VDD DP_OP_655J1_123_1759_n71 DP_OP_655J1_123_1759_n77 DP_OP_655J1_123_1759_n75 DP_OP_655J1_123_1759_n67 DP_OP_655J1_123_1759_n68 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U243 VSS VDD in_data1_dff[120] in_data1_dff[96] in_data1_dff[88] DP_OP_654J1_122_1759_n332 DP_OP_654J1_122_1759_n333 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U242 VSS VDD in_data1_dff[80] in_data1_dff[72] in_data1_dff[64] DP_OP_654J1_122_1759_n330 DP_OP_654J1_122_1759_n331 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U241 VSS VDD in_data1_dff[56] in_data1_dff[48] in_data1_dff[40] DP_OP_654J1_122_1759_n328 DP_OP_654J1_122_1759_n329 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U240 VSS VDD in_data1_dff[32] in_data1_dff[24] in_data1_dff[16] DP_OP_654J1_122_1759_n326 DP_OP_654J1_122_1759_n327 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U239 VSS VDD in_data1_dff[8] in_data1_dff[0] in_data1_dff[4] DP_OP_654J1_122_1759_n324 DP_OP_654J1_122_1759_n325 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U238 VSS VDD in_data1_dff[12] in_data1_dff[20] in_data1_dff[28] DP_OP_654J1_122_1759_n322 DP_OP_654J1_122_1759_n323 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U237 VSS VDD in_data1_dff[36] in_data1_dff[44] in_data1_dff[52] DP_OP_654J1_122_1759_n320 DP_OP_654J1_122_1759_n321 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U236 VSS VDD in_data1_dff[60] in_data1_dff[68] in_data1_dff[76] DP_OP_654J1_122_1759_n318 DP_OP_654J1_122_1759_n319 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U235 VSS VDD in_data1_dff[84] in_data1_dff[124] in_data1_dff[92] DP_OP_654J1_122_1759_n316 DP_OP_654J1_122_1759_n317 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U234 VSS VDD in_data1_dff[100] in_data1_dff[116] in_data1_dff[108] DP_OP_654J1_122_1759_n314 DP_OP_654J1_122_1759_n315 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U232 VSS VDD DP_OP_654J1_122_1759_n317 DP_OP_654J1_122_1759_n311 DP_OP_654J1_122_1759_n319 DP_OP_654J1_122_1759_n312 DP_OP_654J1_122_1759_n313 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U231 VSS VDD DP_OP_654J1_122_1759_n315 DP_OP_654J1_122_1759_n321 DP_OP_654J1_122_1759_n323 DP_OP_654J1_122_1759_n309 DP_OP_654J1_122_1759_n310 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U230 VSS VDD DP_OP_654J1_122_1759_n325 DP_OP_654J1_122_1759_n327 DP_OP_654J1_122_1759_n329 DP_OP_654J1_122_1759_n307 DP_OP_654J1_122_1759_n308 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U228 VSS VDD DP_OP_654J1_122_1759_n331 DP_OP_654J1_122_1759_n333 DP_OP_654J1_122_1759_n304 DP_OP_654J1_122_1759_n305 DP_OP_654J1_122_1759_n306 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U225 VSS VDD in_data1_dff[105] in_data1_dff[97] in_data1_dff[89] DP_OP_654J1_122_1759_n300 DP_OP_654J1_122_1759_n301 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U224 VSS VDD in_data1_dff[81] in_data1_dff[73] in_data1_dff[65] DP_OP_654J1_122_1759_n298 DP_OP_654J1_122_1759_n299 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U223 VSS VDD in_data1_dff[57] in_data1_dff[49] in_data1_dff[41] DP_OP_654J1_122_1759_n296 DP_OP_654J1_122_1759_n297 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U222 VSS VDD in_data1_dff[33] in_data1_dff[25] in_data1_dff[17] DP_OP_654J1_122_1759_n294 DP_OP_654J1_122_1759_n295 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U221 VSS VDD in_data1_dff[9] in_data1_dff[45] in_data1_dff[125] DP_OP_654J1_122_1759_n292 DP_OP_654J1_122_1759_n293 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U220 VSS VDD in_data1_dff[1] in_data1_dff[37] in_data1_dff[5] DP_OP_654J1_122_1759_n290 DP_OP_654J1_122_1759_n291 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U219 VSS VDD in_data1_dff[117] in_data1_dff[61] in_data1_dff[109] DP_OP_654J1_122_1759_n288 DP_OP_654J1_122_1759_n289 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U218 VSS VDD in_data1_dff[13] in_data1_dff[29] in_data1_dff[101] DP_OP_654J1_122_1759_n286 DP_OP_654J1_122_1759_n287 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U217 VSS VDD in_data1_dff[21] in_data1_dff[93] in_data1_dff[53] DP_OP_654J1_122_1759_n284 DP_OP_654J1_122_1759_n285 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U216 VSS VDD in_data1_dff[69] in_data1_dff[85] in_data1_dff[77] DP_OP_654J1_122_1759_n282 DP_OP_654J1_122_1759_n283 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U214 VSS VDD DP_OP_654J1_122_1759_n332 DP_OP_654J1_122_1759_n279 DP_OP_654J1_122_1759_n330 DP_OP_654J1_122_1759_n280 DP_OP_654J1_122_1759_n281 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U212 VSS VDD DP_OP_654J1_122_1759_n328 DP_OP_654J1_122_1759_n316 DP_OP_654J1_122_1759_n276 DP_OP_654J1_122_1759_n277 DP_OP_654J1_122_1759_n278 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U211 VSS VDD DP_OP_654J1_122_1759_n318 DP_OP_654J1_122_1759_n314 DP_OP_654J1_122_1759_n320 DP_OP_654J1_122_1759_n274 DP_OP_654J1_122_1759_n275 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U210 VSS VDD DP_OP_654J1_122_1759_n322 DP_OP_654J1_122_1759_n324 DP_OP_654J1_122_1759_n326 DP_OP_654J1_122_1759_n272 DP_OP_654J1_122_1759_n273 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U209 VSS VDD DP_OP_654J1_122_1759_n293 DP_OP_654J1_122_1759_n283 DP_OP_654J1_122_1759_n295 DP_OP_654J1_122_1759_n270 DP_OP_654J1_122_1759_n271 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U208 VSS VDD DP_OP_654J1_122_1759_n291 DP_OP_654J1_122_1759_n285 DP_OP_654J1_122_1759_n289 DP_OP_654J1_122_1759_n268 DP_OP_654J1_122_1759_n269 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U207 VSS VDD DP_OP_654J1_122_1759_n299 DP_OP_654J1_122_1759_n287 DP_OP_654J1_122_1759_n297 DP_OP_654J1_122_1759_n266 DP_OP_654J1_122_1759_n267 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U205 VSS VDD DP_OP_654J1_122_1759_n312 DP_OP_654J1_122_1759_n281 DP_OP_654J1_122_1759_n263 DP_OP_654J1_122_1759_n264 DP_OP_654J1_122_1759_n265 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U204 VSS VDD DP_OP_654J1_122_1759_n273 DP_OP_654J1_122_1759_n275 DP_OP_654J1_122_1759_n278 DP_OP_654J1_122_1759_n261 DP_OP_654J1_122_1759_n262 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U203 VSS VDD DP_OP_654J1_122_1759_n307 DP_OP_654J1_122_1759_n309 DP_OP_654J1_122_1759_n271 DP_OP_654J1_122_1759_n259 DP_OP_654J1_122_1759_n260 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U201 VSS VDD DP_OP_654J1_122_1759_n267 DP_OP_654J1_122_1759_n269 DP_OP_654J1_122_1759_n256 DP_OP_654J1_122_1759_n257 DP_OP_654J1_122_1759_n258 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U199 VSS VDD DP_OP_654J1_122_1759_n260 DP_OP_654J1_122_1759_n262 DP_OP_654J1_122_1759_n253 DP_OP_654J1_122_1759_n254 DP_OP_654J1_122_1759_n255 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U195 VSS VDD in_data1_dff[106] in_data1_dff[98] in_data1_dff[90] DP_OP_654J1_122_1759_n248 DP_OP_654J1_122_1759_n249 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U194 VSS VDD in_data1_dff[82] in_data1_dff[74] in_data1_dff[66] DP_OP_654J1_122_1759_n246 DP_OP_654J1_122_1759_n247 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U193 VSS VDD in_data1_dff[126] in_data1_dff[22] in_data1_dff[118] DP_OP_654J1_122_1759_n244 DP_OP_654J1_122_1759_n245 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U192 VSS VDD in_data1_dff[58] in_data1_dff[110] in_data1_dff[50] DP_OP_654J1_122_1759_n242 DP_OP_654J1_122_1759_n243 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U191 VSS VDD in_data1_dff[42] in_data1_dff[102] in_data1_dff[94] DP_OP_654J1_122_1759_n240 DP_OP_654J1_122_1759_n241 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U190 VSS VDD in_data1_dff[34] in_data1_dff[6] in_data1_dff[26] DP_OP_654J1_122_1759_n238 DP_OP_654J1_122_1759_n239 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U189 VSS VDD in_data1_dff[18] in_data1_dff[86] in_data1_dff[10] DP_OP_654J1_122_1759_n236 DP_OP_654J1_122_1759_n237 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U188 VSS VDD in_data1_dff[2] in_data1_dff[78] in_data1_dff[14] DP_OP_654J1_122_1759_n234 DP_OP_654J1_122_1759_n235 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U187 VSS VDD in_data1_dff[70] in_data1_dff[38] in_data1_dff[62] DP_OP_654J1_122_1759_n232 DP_OP_654J1_122_1759_n233 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U186 VSS VDD in_data1_dff[30] in_data1_dff[54] in_data1_dff[46] DP_OP_654J1_122_1759_n230 DP_OP_654J1_122_1759_n231 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U184 VSS VDD DP_OP_654J1_122_1759_n300 DP_OP_654J1_122_1759_n227 DP_OP_654J1_122_1759_n298 DP_OP_654J1_122_1759_n228 DP_OP_654J1_122_1759_n229 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U182 VSS VDD DP_OP_654J1_122_1759_n296 DP_OP_654J1_122_1759_n282 DP_OP_654J1_122_1759_n224 DP_OP_654J1_122_1759_n225 DP_OP_654J1_122_1759_n226 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U181 VSS VDD DP_OP_654J1_122_1759_n294 DP_OP_654J1_122_1759_n290 DP_OP_654J1_122_1759_n284 DP_OP_654J1_122_1759_n222 DP_OP_654J1_122_1759_n223 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U180 VSS VDD DP_OP_654J1_122_1759_n292 DP_OP_654J1_122_1759_n286 DP_OP_654J1_122_1759_n288 DP_OP_654J1_122_1759_n220 DP_OP_654J1_122_1759_n221 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U178 VSS VDD DP_OP_654J1_122_1759_n274 DP_OP_654J1_122_1759_n280 DP_OP_654J1_122_1759_n217 DP_OP_654J1_122_1759_n218 DP_OP_654J1_122_1759_n219 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U176 VSS VDD DP_OP_654J1_122_1759_n243 DP_OP_654J1_122_1759_n235 DP_OP_654J1_122_1759_n214 DP_OP_654J1_122_1759_n215 DP_OP_654J1_122_1759_n216 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U175 VSS VDD DP_OP_654J1_122_1759_n247 DP_OP_654J1_122_1759_n237 DP_OP_654J1_122_1759_n249 DP_OP_654J1_122_1759_n212 DP_OP_654J1_122_1759_n213 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U174 VSS VDD DP_OP_654J1_122_1759_n245 DP_OP_654J1_122_1759_n233 DP_OP_654J1_122_1759_n239 DP_OP_654J1_122_1759_n210 DP_OP_654J1_122_1759_n211 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U172 VSS VDD DP_OP_654J1_122_1759_n277 DP_OP_654J1_122_1759_n229 DP_OP_654J1_122_1759_n207 DP_OP_654J1_122_1759_n208 DP_OP_654J1_122_1759_n209 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U171 VSS VDD DP_OP_654J1_122_1759_n223 DP_OP_654J1_122_1759_n221 DP_OP_654J1_122_1759_n226 DP_OP_654J1_122_1759_n205 DP_OP_654J1_122_1759_n206 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U170 VSS VDD DP_OP_654J1_122_1759_n266 DP_OP_654J1_122_1759_n270 DP_OP_654J1_122_1759_n268 DP_OP_654J1_122_1759_n203 DP_OP_654J1_122_1759_n204 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U168 VSS VDD DP_OP_654J1_122_1759_n261 DP_OP_654J1_122_1759_n264 DP_OP_654J1_122_1759_n200 DP_OP_654J1_122_1759_n201 DP_OP_654J1_122_1759_n202 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U166 VSS VDD DP_OP_654J1_122_1759_n213 DP_OP_654J1_122_1759_n211 DP_OP_654J1_122_1759_n197 DP_OP_654J1_122_1759_n198 DP_OP_654J1_122_1759_n199 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U165 VSS VDD DP_OP_654J1_122_1759_n259 DP_OP_654J1_122_1759_n209 DP_OP_654J1_122_1759_n204 DP_OP_654J1_122_1759_n195 DP_OP_654J1_122_1759_n196 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U164 VSS VDD DP_OP_654J1_122_1759_n257 DP_OP_654J1_122_1759_n206 DP_OP_654J1_122_1759_n199 DP_OP_654J1_122_1759_n193 DP_OP_654J1_122_1759_n194 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U163 VSS VDD DP_OP_654J1_122_1759_n254 DP_OP_654J1_122_1759_n202 DP_OP_654J1_122_1759_n196 DP_OP_654J1_122_1759_n191 DP_OP_654J1_122_1759_n192 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U159 VSS VDD in_data1_dff[107] in_data1_dff[99] in_data1_dff[91] DP_OP_654J1_122_1759_n186 DP_OP_654J1_122_1759_n187 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U158 VSS VDD in_data1_dff[83] in_data1_dff[15] in_data1_dff[75] DP_OP_654J1_122_1759_n184 DP_OP_654J1_122_1759_n185 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U157 VSS VDD in_data1_dff[67] in_data1_dff[127] in_data1_dff[59] DP_OP_654J1_122_1759_n182 DP_OP_654J1_122_1759_n183 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U156 VSS VDD in_data1_dff[51] in_data1_dff[31] in_data1_dff[119] DP_OP_654J1_122_1759_n180 DP_OP_654J1_122_1759_n181 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U155 VSS VDD in_data1_dff[111] in_data1_dff[23] in_data1_dff[43] DP_OP_654J1_122_1759_n178 DP_OP_654J1_122_1759_n179 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U154 VSS VDD in_data1_dff[35] in_data1_dff[103] in_data1_dff[27] DP_OP_654J1_122_1759_n176 DP_OP_654J1_122_1759_n177 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U153 VSS VDD in_data1_dff[19] in_data1_dff[95] in_data1_dff[11] DP_OP_654J1_122_1759_n174 DP_OP_654J1_122_1759_n175 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U152 VSS VDD in_data1_dff[3] in_data1_dff[87] in_data1_dff[7] DP_OP_654J1_122_1759_n172 DP_OP_654J1_122_1759_n173 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U151 VSS VDD in_data1_dff[39] in_data1_dff[79] in_data1_dff[47] DP_OP_654J1_122_1759_n170 DP_OP_654J1_122_1759_n171 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U150 VSS VDD in_data1_dff[55] in_data1_dff[71] in_data1_dff[63] DP_OP_654J1_122_1759_n168 DP_OP_654J1_122_1759_n169 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U148 VSS VDD DP_OP_654J1_122_1759_n248 DP_OP_654J1_122_1759_n165 DP_OP_654J1_122_1759_n246 DP_OP_654J1_122_1759_n166 DP_OP_654J1_122_1759_n167 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U146 VSS VDD DP_OP_654J1_122_1759_n244 DP_OP_654J1_122_1759_n230 DP_OP_654J1_122_1759_n162 DP_OP_654J1_122_1759_n163 DP_OP_654J1_122_1759_n164 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U145 VSS VDD DP_OP_654J1_122_1759_n242 DP_OP_654J1_122_1759_n238 DP_OP_654J1_122_1759_n232 DP_OP_654J1_122_1759_n160 DP_OP_654J1_122_1759_n161 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U144 VSS VDD DP_OP_654J1_122_1759_n240 DP_OP_654J1_122_1759_n236 DP_OP_654J1_122_1759_n234 DP_OP_654J1_122_1759_n158 DP_OP_654J1_122_1759_n159 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U142 VSS VDD DP_OP_654J1_122_1759_n222 DP_OP_654J1_122_1759_n228 DP_OP_654J1_122_1759_n155 DP_OP_654J1_122_1759_n156 DP_OP_654J1_122_1759_n157 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U140 VSS VDD DP_OP_654J1_122_1759_n183 DP_OP_654J1_122_1759_n169 DP_OP_654J1_122_1759_n152 DP_OP_654J1_122_1759_n153 DP_OP_654J1_122_1759_n154 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U139 VSS VDD DP_OP_654J1_122_1759_n181 DP_OP_654J1_122_1759_n175 DP_OP_654J1_122_1759_n179 DP_OP_654J1_122_1759_n150 DP_OP_654J1_122_1759_n151 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U138 VSS VDD DP_OP_654J1_122_1759_n185 DP_OP_654J1_122_1759_n187 DP_OP_654J1_122_1759_n177 DP_OP_654J1_122_1759_n148 DP_OP_654J1_122_1759_n149 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U136 VSS VDD DP_OP_654J1_122_1759_n225 DP_OP_654J1_122_1759_n167 DP_OP_654J1_122_1759_n145 DP_OP_654J1_122_1759_n146 DP_OP_654J1_122_1759_n147 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U134 VSS VDD DP_OP_654J1_122_1759_n215 DP_OP_654J1_122_1759_n212 DP_OP_654J1_122_1759_n142 DP_OP_654J1_122_1759_n143 DP_OP_654J1_122_1759_n144 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U133 VSS VDD DP_OP_654J1_122_1759_n161 DP_OP_654J1_122_1759_n210 DP_OP_654J1_122_1759_n164 DP_OP_654J1_122_1759_n140 DP_OP_654J1_122_1759_n141 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U131 VSS VDD DP_OP_654J1_122_1759_n149 DP_OP_654J1_122_1759_n159 DP_OP_654J1_122_1759_n137 DP_OP_654J1_122_1759_n138 DP_OP_654J1_122_1759_n139 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U129 VSS VDD DP_OP_654J1_122_1759_n203 DP_OP_654J1_122_1759_n157 DP_OP_654J1_122_1759_n134 DP_OP_654J1_122_1759_n135 DP_OP_654J1_122_1759_n136 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U127 VSS VDD DP_OP_654J1_122_1759_n205 DP_OP_654J1_122_1759_n147 DP_OP_654J1_122_1759_n131 DP_OP_654J1_122_1759_n132 DP_OP_654J1_122_1759_n133 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U125 VSS VDD DP_OP_654J1_122_1759_n144 DP_OP_654J1_122_1759_n141 DP_OP_654J1_122_1759_n128 DP_OP_654J1_122_1759_n129 DP_OP_654J1_122_1759_n130 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U123 VSS VDD DP_OP_654J1_122_1759_n139 DP_OP_654J1_122_1759_n198 DP_OP_654J1_122_1759_n125 DP_OP_654J1_122_1759_n126 DP_OP_654J1_122_1759_n127 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U122 VSS VDD DP_OP_654J1_122_1759_n133 DP_OP_654J1_122_1759_n136 DP_OP_654J1_122_1759_n193 DP_OP_654J1_122_1759_n123 DP_OP_654J1_122_1759_n124 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U120 VSS VDD DP_OP_654J1_122_1759_n127 DP_OP_654J1_122_1759_n130 DP_OP_654J1_122_1759_n120 DP_OP_654J1_122_1759_n121 DP_OP_654J1_122_1759_n122 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U114 VSS VDD DP_OP_654J1_122_1759_n184 DP_OP_654J1_122_1759_n170 DP_OP_654J1_122_1759_n182 DP_OP_654J1_122_1759_n113 DP_OP_654J1_122_1759_n114 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U113 VSS VDD DP_OP_654J1_122_1759_n180 DP_OP_654J1_122_1759_n176 DP_OP_654J1_122_1759_n168 DP_OP_654J1_122_1759_n111 DP_OP_654J1_122_1759_n112 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U112 VSS VDD DP_OP_654J1_122_1759_n172 DP_OP_654J1_122_1759_n174 DP_OP_654J1_122_1759_n178 DP_OP_654J1_122_1759_n109 DP_OP_654J1_122_1759_n110 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U111 VSS VDD DP_OP_654J1_122_1759_n158 DP_OP_654J1_122_1759_n166 DP_OP_654J1_122_1759_n163 DP_OP_654J1_122_1759_n107 DP_OP_654J1_122_1759_n108 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U110 VSS VDD DP_OP_654J1_122_1759_n117 DP_OP_654J1_122_1759_n160 DP_OP_654J1_122_1759_n148 DP_OP_654J1_122_1759_n105 DP_OP_654J1_122_1759_n106 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U108 VSS VDD DP_OP_654J1_122_1759_n153 DP_OP_654J1_122_1759_n110 DP_OP_654J1_122_1759_n102 DP_OP_654J1_122_1759_n103 DP_OP_654J1_122_1759_n104 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U107 VSS VDD DP_OP_654J1_122_1759_n114 DP_OP_654J1_122_1759_n150 DP_OP_654J1_122_1759_n112 DP_OP_654J1_122_1759_n100 DP_OP_654J1_122_1759_n101 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U106 VSS VDD DP_OP_654J1_122_1759_n108 DP_OP_654J1_122_1759_n146 DP_OP_654J1_122_1759_n140 DP_OP_654J1_122_1759_n98 DP_OP_654J1_122_1759_n99 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U105 VSS VDD DP_OP_654J1_122_1759_n106 DP_OP_654J1_122_1759_n143 DP_OP_654J1_122_1759_n138 DP_OP_654J1_122_1759_n96 DP_OP_654J1_122_1759_n97 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U103 VSS VDD DP_OP_654J1_122_1759_n104 DP_OP_654J1_122_1759_n101 DP_OP_654J1_122_1759_n93 DP_OP_654J1_122_1759_n94 DP_OP_654J1_122_1759_n95 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U102 VSS VDD DP_OP_654J1_122_1759_n99 DP_OP_654J1_122_1759_n132 DP_OP_654J1_122_1759_n129 DP_OP_654J1_122_1759_n91 DP_OP_654J1_122_1759_n92 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U101 VSS VDD DP_OP_654J1_122_1759_n126 DP_OP_654J1_122_1759_n97 DP_OP_654J1_122_1759_n95 DP_OP_654J1_122_1759_n89 DP_OP_654J1_122_1759_n90 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U100 VSS VDD DP_OP_654J1_122_1759_n92 DP_OP_654J1_122_1759_n123 DP_OP_654J1_122_1759_n121 DP_OP_654J1_122_1759_n87 DP_OP_654J1_122_1759_n88 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U98 VSS VDD DP_OP_654J1_122_1759_n109 DP_OP_654J1_122_1759_n116 DP_OP_654J1_122_1759_n113 DP_OP_654J1_122_1759_n84 DP_OP_654J1_122_1759_n85 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U96 VSS VDD DP_OP_654J1_122_1759_n107 DP_OP_654J1_122_1759_n105 DP_OP_654J1_122_1759_n81 DP_OP_654J1_122_1759_n82 DP_OP_654J1_122_1759_n83 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U95 VSS VDD DP_OP_654J1_122_1759_n100 DP_OP_654J1_122_1759_n85 DP_OP_654J1_122_1759_n103 DP_OP_654J1_122_1759_n79 DP_OP_654J1_122_1759_n80 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U94 VSS VDD DP_OP_654J1_122_1759_n83 DP_OP_654J1_122_1759_n98 DP_OP_654J1_122_1759_n96 DP_OP_654J1_122_1759_n77 DP_OP_654J1_122_1759_n78 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U92 VSS VDD DP_OP_654J1_122_1759_n94 DP_OP_654J1_122_1759_n80 DP_OP_654J1_122_1759_n74 DP_OP_654J1_122_1759_n75 DP_OP_654J1_122_1759_n76 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U91 VSS VDD DP_OP_654J1_122_1759_n89 DP_OP_654J1_122_1759_n78 DP_OP_654J1_122_1759_n76 DP_OP_654J1_122_1759_n72 DP_OP_654J1_122_1759_n73 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U89 VSS VDD DP_OP_654J1_122_1759_n82 DP_OP_654J1_122_1759_n79 DP_OP_654J1_122_1759_n69 DP_OP_654J1_122_1759_n70 DP_OP_654J1_122_1759_n71 FAx1_ASAP7_75t_R
XDP_OP_654J1_122_1759_U88 VSS VDD DP_OP_654J1_122_1759_n71 DP_OP_654J1_122_1759_n77 DP_OP_654J1_122_1759_n75 DP_OP_654J1_122_1759_n67 DP_OP_654J1_122_1759_n68 FAx1_ASAP7_75t_R
XU1840 VSS VDD DP_OP_654J1_122_1759_n258 n1091 n1020 A0 n1092 FAx1_ASAP7_75t_R
XU1845 VSS VDD DP_OP_655J1_123_1759_n258 n1098 n1022 A2 n1099 FAx1_ASAP7_75t_R
XU1850 VSS VDD DP_OP_657J1_125_1759_n258 n1112 n1017 A4 n1113 FAx1_ASAP7_75t_R
XU1855 VSS VDD DP_OP_656J1_124_1759_n258 n1105 n1024 A6 n1106 FAx1_ASAP7_75t_R
XU1860 VSS VDD n1141 DP_OP_654J1_122_1759_n194 n1003 A8 n1138 FAx1_ASAP7_75t_R
XU1867 VSS VDD n1132 DP_OP_655J1_123_1759_n194 n1005 A10 n1129 FAx1_ASAP7_75t_R
XU1874 VSS VDD n1123 DP_OP_656J1_124_1759_n194 n994 A12 n1120 FAx1_ASAP7_75t_R
XU1881 VSS VDD n1149 DP_OP_657J1_125_1759_n194 n996 A14 n1146 FAx1_ASAP7_75t_R
XU1889 VSS VDD DP_OP_656J1_124_1759_n122 DP_OP_656J1_124_1759_n124 n935 A17 n1161 FAx1_ASAP7_75t_R
XU1894 VSS VDD DP_OP_655J1_123_1759_n122 DP_OP_655J1_123_1759_n124 n936 A20 n1168 FAx1_ASAP7_75t_R
XU1900 VSS VDD DP_OP_654J1_122_1759_n122 DP_OP_654J1_122_1759_n124 n933 A23 n1175 FAx1_ASAP7_75t_R
XU1906 VSS VDD DP_OP_657J1_125_1759_n122 DP_OP_657J1_125_1759_n124 n934 A26 n1154 FAx1_ASAP7_75t_R
XU1911 VSS VDD n1186 DP_OP_657J1_125_1759_n88 n1000 A28 n1184 FAx1_ASAP7_75t_R
XU1918 VSS VDD n1203 DP_OP_656J1_124_1759_n88 n992 A30 n1201 FAx1_ASAP7_75t_R
XU1925 VSS VDD n1212 DP_OP_655J1_123_1759_n88 n998 A32 n1210 FAx1_ASAP7_75t_R
XU1932 VSS VDD n1194 DP_OP_654J1_122_1759_n88 n990 A34 n1192 FAx1_ASAP7_75t_R
XU1940 VSS VDD n1217 DP_OP_657J1_125_1759_n87 DP_OP_657J1_125_1759_n73 A37 n1218 FAx1_ASAP7_75t_R
XU1945 VSS VDD n1225 DP_OP_654J1_122_1759_n87 DP_OP_654J1_122_1759_n73 A40 n1226 FAx1_ASAP7_75t_R
XU1950 VSS VDD n1241 DP_OP_656J1_124_1759_n87 DP_OP_656J1_124_1759_n73 A43 n1242 FAx1_ASAP7_75t_R
XU1955 VSS VDD n1233 DP_OP_655J1_123_1759_n87 DP_OP_655J1_123_1759_n73 A46 n1234 FAx1_ASAP7_75t_R
XU1958 VSS VDD DP_OP_657J1_125_1759_n72 DP_OP_657J1_125_1759_n68 n917 A48 n1251 FAx1_ASAP7_75t_R
XU1964 VSS VDD DP_OP_654J1_122_1759_n72 DP_OP_654J1_122_1759_n68 n916 A50 n1260 FAx1_ASAP7_75t_R
XU1970 VSS VDD DP_OP_655J1_123_1759_n72 DP_OP_655J1_123_1759_n68 n914 A52 n1269 FAx1_ASAP7_75t_R
XU1976 VSS VDD DP_OP_656J1_124_1759_n72 DP_OP_656J1_124_1759_n68 n915 A54 n1278 FAx1_ASAP7_75t_R
XU1985 VSS VDD DP_OP_657J1_125_1759_n70 n1053 n1294 A57 n1295 FAx1_ASAP7_75t_R
XU1991 VSS VDD DP_OP_654J1_122_1759_n70 n1054 n1286 A60 n1287 FAx1_ASAP7_75t_R
XU1997 VSS VDD DP_OP_655J1_123_1759_n70 n1055 n1302 A63 n1303 FAx1_ASAP7_75t_R
XU2003 VSS VDD DP_OP_656J1_124_1759_n70 n1056 n1310 A66 n1311 FAx1_ASAP7_75t_R
XU1841 VSS VDD n1075 n1092 A1 n1076 HAxp5_ASAP7_75t_R
XU1846 VSS VDD n1079 n1099 A3 n1080 HAxp5_ASAP7_75t_R
XU1851 VSS VDD n1083 n1113 A5 n1084 HAxp5_ASAP7_75t_R
XU1856 VSS VDD n1087 n1106 A7 n1088 HAxp5_ASAP7_75t_R
XU1862 VSS VDD n1139 n1137 A9 n1093 HAxp5_ASAP7_75t_R
XU1869 VSS VDD n1130 n1128 A11 n1100 HAxp5_ASAP7_75t_R
XU1876 VSS VDD n1121 n1119 A13 n1107 HAxp5_ASAP7_75t_R
XU1883 VSS VDD n1147 n956 A15 n1114 HAxp5_ASAP7_75t_R
XU1887 VSS VDD n187 n1162 A16 n1122 HAxp5_ASAP7_75t_R
XU1890 VSS VDD n1124 n1161 A18 n1125 HAxp5_ASAP7_75t_R
XU1892 VSS VDD n213 n1169 A19 n1131 HAxp5_ASAP7_75t_R
XU1895 VSS VDD n1133 n1168 A21 n1134 HAxp5_ASAP7_75t_R
XU1898 VSS VDD n239 n1176 A22 n1140 HAxp5_ASAP7_75t_R
XU1901 VSS VDD n1142 n1175 A24 n1143 HAxp5_ASAP7_75t_R
XU1904 VSS VDD n265 n1155 A25 n1148 HAxp5_ASAP7_75t_R
XU1907 VSS VDD n1150 n1154 A27 n1151 HAxp5_ASAP7_75t_R
XU1913 VSS VDD n1183 n1182 A29 n1156 HAxp5_ASAP7_75t_R
XU1920 VSS VDD n1200 n1199 A31 n1163 HAxp5_ASAP7_75t_R
XU1927 VSS VDD n1209 n1208 A33 n1170 HAxp5_ASAP7_75t_R
XU1934 VSS VDD n1191 n957 A35 n1177 HAxp5_ASAP7_75t_R
XU1938 VSS VDD n269 n1219 A36 n1185 HAxp5_ASAP7_75t_R
XU1941 VSS VDD n1187 n1218 A38 n1188 HAxp5_ASAP7_75t_R
XU1943 VSS VDD n243 n1227 A39 n1193 HAxp5_ASAP7_75t_R
XU1946 VSS VDD n1195 n1226 A41 n1196 HAxp5_ASAP7_75t_R
XU1948 VSS VDD n191 n1243 A42 n1202 HAxp5_ASAP7_75t_R
XU1951 VSS VDD n1204 n1242 A44 n1205 HAxp5_ASAP7_75t_R
XU1953 VSS VDD n217 n1235 A45 n1211 HAxp5_ASAP7_75t_R
XU1956 VSS VDD n1213 n1234 A47 n1214 HAxp5_ASAP7_75t_R
XU1960 VSS VDD n1250 n1042 A49 n1220 HAxp5_ASAP7_75t_R
XU1966 VSS VDD n1259 n1043 A51 n1228 HAxp5_ASAP7_75t_R
XU1972 VSS VDD n1268 n1267 A53 n1236 HAxp5_ASAP7_75t_R
XU1978 VSS VDD n1277 n1044 A55 n1244 HAxp5_ASAP7_75t_R
XU1982 VSS VDD n273 n1296 A56 n1252 HAxp5_ASAP7_75t_R
XU1986 VSS VDD n1254 n1295 A58 n1255 HAxp5_ASAP7_75t_R
XU1988 VSS VDD n247 n1288 A59 n1261 HAxp5_ASAP7_75t_R
XU1992 VSS VDD n1263 n1287 A61 n1264 HAxp5_ASAP7_75t_R
XU1994 VSS VDD n221 n1304 A62 n1270 HAxp5_ASAP7_75t_R
XU1998 VSS VDD n1272 n1303 A64 n1273 HAxp5_ASAP7_75t_R
XU2000 VSS VDD n195 n1312 A65 n1279 HAxp5_ASAP7_75t_R
XU2004 VSS VDD n1281 n1311 A67 n1282 HAxp5_ASAP7_75t_R
XU2035 VSS VDD n1337 n1338 A68 n1339 HAxp5_ASAP7_75t_R
XU2039 VSS VDD n1345 n955 A69 n1346 HAxp5_ASAP7_75t_R
XU2043 VSS VDD n1352 n1353 A70 n1354 HAxp5_ASAP7_75t_R
XU2047 VSS VDD n1360 n1361 A71 n1362 HAxp5_ASAP7_75t_R
XU2062 VSS VDD n1384 n205 A72 n1385 HAxp5_ASAP7_75t_R
XU2088 VSS VDD n1388 n231 A73 n1389 HAxp5_ASAP7_75t_R
XU2114 VSS VDD n1392 n257 A74 n1393 HAxp5_ASAP7_75t_R
XU2140 VSS VDD n1396 n283 A75 n1397 HAxp5_ASAP7_75t_R
XU2168 VSS VDD in_data1_dff[123] in_data1_dff[115] A76 DP_OP_654J1_122_1759_n162 HAxp5_ASAP7_75t_R
XU2169 VSS VDD in_data1_dff[122] in_data1_dff[114] A77 DP_OP_654J1_122_1759_n224 HAxp5_ASAP7_75t_R
XU2170 VSS VDD in_data1_dff[121] in_data1_dff[113] A78 DP_OP_654J1_122_1759_n276 HAxp5_ASAP7_75t_R
XU2171 VSS VDD in_data1_dff[112] in_data1_dff[104] A79 DP_OP_654J1_122_1759_n311 HAxp5_ASAP7_75t_R
XU2174 VSS VDD in_data2_dff[123] in_data2_dff[115] A80 DP_OP_655J1_123_1759_n162 HAxp5_ASAP7_75t_R
XU2175 VSS VDD in_data2_dff[122] in_data2_dff[114] A81 DP_OP_655J1_123_1759_n224 HAxp5_ASAP7_75t_R
XU2176 VSS VDD in_data2_dff[121] in_data2_dff[113] A82 DP_OP_655J1_123_1759_n276 HAxp5_ASAP7_75t_R
XU2177 VSS VDD in_data2_dff[112] in_data2_dff[104] A83 DP_OP_655J1_123_1759_n311 HAxp5_ASAP7_75t_R
XU2180 VSS VDD in_data3_dff[123] in_data3_dff[115] A84 DP_OP_656J1_124_1759_n162 HAxp5_ASAP7_75t_R
XU2181 VSS VDD in_data3_dff[122] in_data3_dff[114] A85 DP_OP_656J1_124_1759_n224 HAxp5_ASAP7_75t_R
XU2182 VSS VDD in_data3_dff[121] in_data3_dff[113] A86 DP_OP_656J1_124_1759_n276 HAxp5_ASAP7_75t_R
XU2183 VSS VDD in_data3_dff[112] in_data3_dff[104] A87 DP_OP_656J1_124_1759_n311 HAxp5_ASAP7_75t_R
XU2186 VSS VDD in_data4_dff[123] in_data4_dff[115] A88 DP_OP_657J1_125_1759_n162 HAxp5_ASAP7_75t_R
XU2187 VSS VDD in_data4_dff[122] in_data4_dff[114] A89 DP_OP_657J1_125_1759_n224 HAxp5_ASAP7_75t_R
XU2188 VSS VDD in_data4_dff[121] in_data4_dff[113] A90 DP_OP_657J1_125_1759_n276 HAxp5_ASAP7_75t_R
XU2189 VSS VDD in_data4_dff[112] in_data4_dff[104] A91 DP_OP_657J1_125_1759_n311 HAxp5_ASAP7_75t_R
XU2242 VSS VDD n289 n861 A92 n290 HAxp5_ASAP7_75t_R
XU2244 VSS VDD n287 n1405 A93 n288 HAxp5_ASAP7_75t_R
XU2064 VSS VDD DP_OP_656J1_124_1759_n91 DP_OP_656J1_124_1759_n74 INVx1_ASAP7_75t_R
XU2065 VSS VDD DP_OP_656J1_124_1759_n191 DP_OP_656J1_124_1759_n120 INVx1_ASAP7_75t_R
XU2066 VSS VDD DP_OP_656J1_124_1759_n305 DP_OP_656J1_124_1759_n253 INVx1_ASAP7_75t_R
XU2067 VSS VDD DP_OP_656J1_124_1759_n313 DP_OP_656J1_124_1759_n304 INVx1_ASAP7_75t_R
XU2068 VSS VDD DP_OP_656J1_124_1759_n201 DP_OP_656J1_124_1759_n128 INVx1_ASAP7_75t_R
XU2069 VSS VDD DP_OP_656J1_124_1759_n216 DP_OP_656J1_124_1759_n200 INVx1_ASAP7_75t_R
XU2070 VSS VDD DP_OP_656J1_124_1759_n265 DP_OP_656J1_124_1759_n256 INVx1_ASAP7_75t_R
XU2071 VSS VDD DP_OP_656J1_124_1759_n301 DP_OP_656J1_124_1759_n263 INVx1_ASAP7_75t_R
XU2072 VSS VDD DP_OP_656J1_124_1759_n171 DP_OP_656J1_124_1759_n145 INVx1_ASAP7_75t_R
XU2073 VSS VDD DP_OP_656J1_124_1759_n154 DP_OP_656J1_124_1759_n131 INVx1_ASAP7_75t_R
XU2074 VSS VDD DP_OP_656J1_124_1759_n135 DP_OP_656J1_124_1759_n93 INVx1_ASAP7_75t_R
XU2075 VSS VDD DP_OP_656J1_124_1759_n151 DP_OP_656J1_124_1759_n134 INVx1_ASAP7_75t_R
XU2076 VSS VDD DP_OP_656J1_124_1759_n218 DP_OP_656J1_124_1759_n142 INVx1_ASAP7_75t_R
XU2077 VSS VDD DP_OP_656J1_124_1759_n272 DP_OP_656J1_124_1759_n214 INVx1_ASAP7_75t_R
XU2078 VSS VDD DP_OP_656J1_124_1759_n195 DP_OP_656J1_124_1759_n125 INVx1_ASAP7_75t_R
XU2079 VSS VDD DP_OP_656J1_124_1759_n219 DP_OP_656J1_124_1759_n197 INVx1_ASAP7_75t_R
XU2080 VSS VDD DP_OP_656J1_124_1759_n231 DP_OP_656J1_124_1759_n217 INVx1_ASAP7_75t_R
XU2081 VSS VDD DP_OP_656J1_124_1759_n208 DP_OP_656J1_124_1759_n137 INVx1_ASAP7_75t_R
XU2082 VSS VDD DP_OP_656J1_124_1759_n241 DP_OP_656J1_124_1759_n207 INVx1_ASAP7_75t_R
XU2083 VSS VDD DP_OP_656J1_124_1759_n156 DP_OP_656J1_124_1759_n102 INVx1_ASAP7_75t_R
XU2084 VSS VDD DP_OP_656J1_124_1759_n173 DP_OP_656J1_124_1759_n155 INVx1_ASAP7_75t_R
XU2085 VSS VDD DP_OP_656J1_124_1759_n220 DP_OP_656J1_124_1759_n152 INVx1_ASAP7_75t_R
XU2086 VSS VDD DP_OP_656J1_124_1759_n84 DP_OP_656J1_124_1759_n69 INVx1_ASAP7_75t_R
XU2087 VSS VDD DP_OP_656J1_124_1759_n111 DP_OP_656J1_124_1759_n81 INVx1_ASAP7_75t_R
XU2090 VSS VDD DP_OP_655J1_123_1759_n91 DP_OP_655J1_123_1759_n74 INVx1_ASAP7_75t_R
XU2091 VSS VDD DP_OP_655J1_123_1759_n191 DP_OP_655J1_123_1759_n120 INVx1_ASAP7_75t_R
XU2092 VSS VDD DP_OP_655J1_123_1759_n305 DP_OP_655J1_123_1759_n253 INVx1_ASAP7_75t_R
XU2093 VSS VDD DP_OP_655J1_123_1759_n313 DP_OP_655J1_123_1759_n304 INVx1_ASAP7_75t_R
XU2094 VSS VDD DP_OP_655J1_123_1759_n201 DP_OP_655J1_123_1759_n128 INVx1_ASAP7_75t_R
XU2095 VSS VDD DP_OP_655J1_123_1759_n216 DP_OP_655J1_123_1759_n200 INVx1_ASAP7_75t_R
XU2096 VSS VDD DP_OP_655J1_123_1759_n265 DP_OP_655J1_123_1759_n256 INVx1_ASAP7_75t_R
XU2097 VSS VDD DP_OP_655J1_123_1759_n301 DP_OP_655J1_123_1759_n263 INVx1_ASAP7_75t_R
XU2098 VSS VDD DP_OP_655J1_123_1759_n171 DP_OP_655J1_123_1759_n145 INVx1_ASAP7_75t_R
XU2099 VSS VDD DP_OP_655J1_123_1759_n154 DP_OP_655J1_123_1759_n131 INVx1_ASAP7_75t_R
XU2100 VSS VDD DP_OP_655J1_123_1759_n135 DP_OP_655J1_123_1759_n93 INVx1_ASAP7_75t_R
XU2101 VSS VDD DP_OP_655J1_123_1759_n151 DP_OP_655J1_123_1759_n134 INVx1_ASAP7_75t_R
XU2102 VSS VDD DP_OP_655J1_123_1759_n218 DP_OP_655J1_123_1759_n142 INVx1_ASAP7_75t_R
XU2103 VSS VDD DP_OP_655J1_123_1759_n272 DP_OP_655J1_123_1759_n214 INVx1_ASAP7_75t_R
XU2104 VSS VDD DP_OP_655J1_123_1759_n195 DP_OP_655J1_123_1759_n125 INVx1_ASAP7_75t_R
XU2105 VSS VDD DP_OP_655J1_123_1759_n219 DP_OP_655J1_123_1759_n197 INVx1_ASAP7_75t_R
XU2106 VSS VDD DP_OP_655J1_123_1759_n231 DP_OP_655J1_123_1759_n217 INVx1_ASAP7_75t_R
XU2107 VSS VDD DP_OP_655J1_123_1759_n208 DP_OP_655J1_123_1759_n137 INVx1_ASAP7_75t_R
XU2108 VSS VDD DP_OP_655J1_123_1759_n241 DP_OP_655J1_123_1759_n207 INVx1_ASAP7_75t_R
XU2109 VSS VDD DP_OP_655J1_123_1759_n156 DP_OP_655J1_123_1759_n102 INVx1_ASAP7_75t_R
XU2110 VSS VDD DP_OP_655J1_123_1759_n173 DP_OP_655J1_123_1759_n155 INVx1_ASAP7_75t_R
XU2111 VSS VDD DP_OP_655J1_123_1759_n220 DP_OP_655J1_123_1759_n152 INVx1_ASAP7_75t_R
XU2112 VSS VDD DP_OP_655J1_123_1759_n84 DP_OP_655J1_123_1759_n69 INVx1_ASAP7_75t_R
XU2113 VSS VDD DP_OP_655J1_123_1759_n111 DP_OP_655J1_123_1759_n81 INVx1_ASAP7_75t_R
XU2116 VSS VDD DP_OP_654J1_122_1759_n91 DP_OP_654J1_122_1759_n74 INVx1_ASAP7_75t_R
XU2117 VSS VDD DP_OP_654J1_122_1759_n191 DP_OP_654J1_122_1759_n120 INVx1_ASAP7_75t_R
XU2118 VSS VDD DP_OP_654J1_122_1759_n305 DP_OP_654J1_122_1759_n253 INVx1_ASAP7_75t_R
XU2119 VSS VDD DP_OP_654J1_122_1759_n313 DP_OP_654J1_122_1759_n304 INVx1_ASAP7_75t_R
XU2120 VSS VDD DP_OP_654J1_122_1759_n201 DP_OP_654J1_122_1759_n128 INVx1_ASAP7_75t_R
XU2121 VSS VDD DP_OP_654J1_122_1759_n216 DP_OP_654J1_122_1759_n200 INVx1_ASAP7_75t_R
XU2122 VSS VDD DP_OP_654J1_122_1759_n265 DP_OP_654J1_122_1759_n256 INVx1_ASAP7_75t_R
XU2123 VSS VDD DP_OP_654J1_122_1759_n301 DP_OP_654J1_122_1759_n263 INVx1_ASAP7_75t_R
XU2124 VSS VDD DP_OP_654J1_122_1759_n171 DP_OP_654J1_122_1759_n145 INVx1_ASAP7_75t_R
XU2125 VSS VDD DP_OP_654J1_122_1759_n154 DP_OP_654J1_122_1759_n131 INVx1_ASAP7_75t_R
XU2126 VSS VDD DP_OP_654J1_122_1759_n135 DP_OP_654J1_122_1759_n93 INVx1_ASAP7_75t_R
XU2127 VSS VDD DP_OP_654J1_122_1759_n151 DP_OP_654J1_122_1759_n134 INVx1_ASAP7_75t_R
XU2128 VSS VDD DP_OP_654J1_122_1759_n218 DP_OP_654J1_122_1759_n142 INVx1_ASAP7_75t_R
XU2129 VSS VDD DP_OP_654J1_122_1759_n272 DP_OP_654J1_122_1759_n214 INVx1_ASAP7_75t_R
XU2130 VSS VDD DP_OP_654J1_122_1759_n195 DP_OP_654J1_122_1759_n125 INVx1_ASAP7_75t_R
XU2131 VSS VDD DP_OP_654J1_122_1759_n219 DP_OP_654J1_122_1759_n197 INVx1_ASAP7_75t_R
XU2132 VSS VDD DP_OP_654J1_122_1759_n231 DP_OP_654J1_122_1759_n217 INVx1_ASAP7_75t_R
XU2133 VSS VDD DP_OP_654J1_122_1759_n208 DP_OP_654J1_122_1759_n137 INVx1_ASAP7_75t_R
XU2134 VSS VDD DP_OP_654J1_122_1759_n241 DP_OP_654J1_122_1759_n207 INVx1_ASAP7_75t_R
XU2135 VSS VDD DP_OP_654J1_122_1759_n156 DP_OP_654J1_122_1759_n102 INVx1_ASAP7_75t_R
XU2136 VSS VDD DP_OP_654J1_122_1759_n173 DP_OP_654J1_122_1759_n155 INVx1_ASAP7_75t_R
XU2137 VSS VDD DP_OP_654J1_122_1759_n220 DP_OP_654J1_122_1759_n152 INVx1_ASAP7_75t_R
XU2138 VSS VDD DP_OP_654J1_122_1759_n84 DP_OP_654J1_122_1759_n69 INVx1_ASAP7_75t_R
XU2139 VSS VDD DP_OP_654J1_122_1759_n111 DP_OP_654J1_122_1759_n81 INVx1_ASAP7_75t_R
XU2142 VSS VDD DP_OP_657J1_125_1759_n91 DP_OP_657J1_125_1759_n74 INVx1_ASAP7_75t_R
XU2143 VSS VDD DP_OP_657J1_125_1759_n191 DP_OP_657J1_125_1759_n120 INVx1_ASAP7_75t_R
XU2144 VSS VDD DP_OP_657J1_125_1759_n305 DP_OP_657J1_125_1759_n253 INVx1_ASAP7_75t_R
XU2145 VSS VDD DP_OP_657J1_125_1759_n313 DP_OP_657J1_125_1759_n304 INVx1_ASAP7_75t_R
XU2146 VSS VDD DP_OP_657J1_125_1759_n201 DP_OP_657J1_125_1759_n128 INVx1_ASAP7_75t_R
XU2147 VSS VDD DP_OP_657J1_125_1759_n216 DP_OP_657J1_125_1759_n200 INVx1_ASAP7_75t_R
XU2148 VSS VDD DP_OP_657J1_125_1759_n265 DP_OP_657J1_125_1759_n256 INVx1_ASAP7_75t_R
XU2149 VSS VDD DP_OP_657J1_125_1759_n301 DP_OP_657J1_125_1759_n263 INVx1_ASAP7_75t_R
XU2150 VSS VDD DP_OP_657J1_125_1759_n171 DP_OP_657J1_125_1759_n145 INVx1_ASAP7_75t_R
XU2151 VSS VDD DP_OP_657J1_125_1759_n154 DP_OP_657J1_125_1759_n131 INVx1_ASAP7_75t_R
XU2152 VSS VDD DP_OP_657J1_125_1759_n135 DP_OP_657J1_125_1759_n93 INVx1_ASAP7_75t_R
XU2153 VSS VDD DP_OP_657J1_125_1759_n151 DP_OP_657J1_125_1759_n134 INVx1_ASAP7_75t_R
XU2154 VSS VDD DP_OP_657J1_125_1759_n218 DP_OP_657J1_125_1759_n142 INVx1_ASAP7_75t_R
XU2155 VSS VDD DP_OP_657J1_125_1759_n272 DP_OP_657J1_125_1759_n214 INVx1_ASAP7_75t_R
XU2156 VSS VDD DP_OP_657J1_125_1759_n195 DP_OP_657J1_125_1759_n125 INVx1_ASAP7_75t_R
XU2157 VSS VDD DP_OP_657J1_125_1759_n219 DP_OP_657J1_125_1759_n197 INVx1_ASAP7_75t_R
XU2158 VSS VDD DP_OP_657J1_125_1759_n231 DP_OP_657J1_125_1759_n217 INVx1_ASAP7_75t_R
XU2159 VSS VDD DP_OP_657J1_125_1759_n208 DP_OP_657J1_125_1759_n137 INVx1_ASAP7_75t_R
XU2160 VSS VDD DP_OP_657J1_125_1759_n241 DP_OP_657J1_125_1759_n207 INVx1_ASAP7_75t_R
XU2161 VSS VDD DP_OP_657J1_125_1759_n156 DP_OP_657J1_125_1759_n102 INVx1_ASAP7_75t_R
XU2162 VSS VDD DP_OP_657J1_125_1759_n173 DP_OP_657J1_125_1759_n155 INVx1_ASAP7_75t_R
XU2163 VSS VDD DP_OP_657J1_125_1759_n220 DP_OP_657J1_125_1759_n152 INVx1_ASAP7_75t_R
XU2164 VSS VDD DP_OP_657J1_125_1759_n84 DP_OP_657J1_125_1759_n69 INVx1_ASAP7_75t_R
XU2165 VSS VDD DP_OP_657J1_125_1759_n111 DP_OP_657J1_125_1759_n81 INVx1_ASAP7_75t_R
XU916 VSS VDD n989 n990 INVx2_ASAP7_75t_R
XU917 VSS VDD n997 n998 INVx2_ASAP7_75t_R
XU918 VSS VDD n999 n1000 INVx2_ASAP7_75t_R
XU919 VSS VDD n991 n992 INVx2_ASAP7_75t_R
XU920 VSS VDD DP_OP_656J1_124_1759_n90 n991 INVx2_ASAP7_75t_R
XU921 VSS VDD DP_OP_654J1_122_1759_n90 n989 INVx2_ASAP7_75t_R
XU922 VSS VDD DP_OP_655J1_123_1759_n90 n997 INVx2_ASAP7_75t_R
XU923 VSS VDD DP_OP_657J1_125_1759_n90 n999 INVx2_ASAP7_75t_R
XU924 VSS VDD n1004 n1005 INVx2_ASAP7_75t_R
XU925 VSS VDD n993 n994 INVx2_ASAP7_75t_R
XU926 VSS VDD n1002 n1003 INVx2_ASAP7_75t_R
XU927 VSS VDD n995 n996 INVx2_ASAP7_75t_R
XU928 VSS VDD n1021 n1022 INVx2_ASAP7_75t_R
XU929 VSS VDD n1019 n1020 INVx2_ASAP7_75t_R
XU930 VSS VDD n1023 n1024 INVx2_ASAP7_75t_R
XU931 VSS VDD n1016 n1017 INVx2_ASAP7_75t_R
XU932 VSS VDD DP_OP_657J1_125_1759_n192 n995 INVx2_ASAP7_75t_R
XU933 VSS VDD DP_OP_655J1_123_1759_n192 n1004 INVx2_ASAP7_75t_R
XU934 VSS VDD DP_OP_656J1_124_1759_n192 n993 INVx2_ASAP7_75t_R
XU935 VSS VDD DP_OP_654J1_122_1759_n192 n1002 INVx2_ASAP7_75t_R
XU936 VSS VDD DP_OP_657J1_125_1759_n255 n1016 INVx2_ASAP7_75t_R
XU937 VSS VDD DP_OP_655J1_123_1759_n255 n1021 INVx2_ASAP7_75t_R
XU938 VSS VDD DP_OP_654J1_122_1759_n255 n1019 INVx2_ASAP7_75t_R
XU939 VSS VDD DP_OP_656J1_124_1759_n255 n1023 INVx2_ASAP7_75t_R
XU946 VSS VDD n1046 n1327 INVx2_ASAP7_75t_R
XU947 VSS VDD n1048 n1322 INVx2_ASAP7_75t_R
XU948 VSS VDD n1045 n1332 INVx2_ASAP7_75t_R
XU949 VSS VDD n1047 n1317 INVx2_ASAP7_75t_R
XU1082 VSS VDD n1031 n955 INVx4_ASAP7_75t_R
XU1136 VSS VDD n1027 n956 INVx4_ASAP7_75t_R
XU1137 VSS VDD n1029 n957 INVx4_ASAP7_75t_R
XU1204 VSS VDD n1258 n1043 INVx4_ASAP7_75t_R
XU1205 VSS VDD n1249 n1042 INVx4_ASAP7_75t_R
XU1206 VSS VDD n1276 n1044 INVx4_ASAP7_75t_R
XU1207 VSS VDD n1035 n1338 INVx4_ASAP7_75t_R
XU1209 VSS VDD n1028 n1361 INVx4_ASAP7_75t_R
XU1211 VSS VDD n1025 n1353 INVx4_ASAP7_75t_R
XU1213 VSS VDD n1030 n1137 INVx4_ASAP7_75t_R
XU1215 VSS VDD n1034 n1128 INVx4_ASAP7_75t_R
XU1217 VSS VDD n1037 n1119 INVx4_ASAP7_75t_R
XU1219 VSS VDD n1033 n1208 INVx4_ASAP7_75t_R
XU1221 VSS VDD n1032 n1267 INVx4_ASAP7_75t_R
XU1223 VSS VDD n1036 n1199 INVx4_ASAP7_75t_R
XU1225 VSS VDD n1026 n1182 INVx4_ASAP7_75t_R
XU907 VSS VDD n1057 n860 INVx5_ASAP7_75t_R
XU941 VSS VDD n1057 n861 INVx8_ASAP7_75t_R
XU1083 VSS VDD rst_n n864 INVx8_ASAP7_75t_R
XU1084 VSS VDD rst_n n865 INVx8_ASAP7_75t_R
XU1085 VSS VDD rst_n n866 INVx8_ASAP7_75t_R
XU1086 VSS VDD rst_n n867 INVx8_ASAP7_75t_R
XU1087 VSS VDD rst_n n868 INVx8_ASAP7_75t_R
XU1088 VSS VDD rst_n n869 INVx8_ASAP7_75t_R
XU1089 VSS VDD rst_n n870 INVx8_ASAP7_75t_R
XU1090 VSS VDD rst_n n871 INVx8_ASAP7_75t_R
XU1091 VSS VDD rst_n n872 INVx8_ASAP7_75t_R
XU1092 VSS VDD rst_n n873 INVx8_ASAP7_75t_R
XU1093 VSS VDD rst_n n874 INVx8_ASAP7_75t_R
XU1094 VSS VDD rst_n n875 INVx8_ASAP7_75t_R
XU1095 VSS VDD rst_n n876 INVx8_ASAP7_75t_R
XU1096 VSS VDD rst_n n877 INVx8_ASAP7_75t_R
XU1097 VSS VDD rst_n n878 INVx8_ASAP7_75t_R
XU1098 VSS VDD rst_n n879 INVx8_ASAP7_75t_R
XU1099 VSS VDD rst_n n880 INVx8_ASAP7_75t_R
XU1100 VSS VDD rst_n n881 INVx8_ASAP7_75t_R
XU1101 VSS VDD rst_n n882 INVx8_ASAP7_75t_R
XU1102 VSS VDD rst_n n883 INVx8_ASAP7_75t_R
XU1103 VSS VDD rst_n n884 INVx8_ASAP7_75t_R
XU1104 VSS VDD rst_n n885 INVx8_ASAP7_75t_R
XU1105 VSS VDD rst_n n886 INVx8_ASAP7_75t_R
XU1106 VSS VDD rst_n n887 INVx8_ASAP7_75t_R
XU1107 VSS VDD rst_n n888 INVx8_ASAP7_75t_R
XU1108 VSS VDD rst_n n889 INVx8_ASAP7_75t_R
XU1109 VSS VDD rst_n n890 INVx8_ASAP7_75t_R
XU1110 VSS VDD rst_n n891 INVx8_ASAP7_75t_R
XU1111 VSS VDD rst_n n892 INVx8_ASAP7_75t_R
XU1112 VSS VDD rst_n n893 INVx8_ASAP7_75t_R
XU1113 VSS VDD rst_n n894 INVx8_ASAP7_75t_R
XU1114 VSS VDD rst_n n895 INVx8_ASAP7_75t_R
XU1115 VSS VDD rst_n n896 INVx8_ASAP7_75t_R
XU1116 VSS VDD rst_n n897 INVx8_ASAP7_75t_R
XU1117 VSS VDD rst_n n898 INVx8_ASAP7_75t_R
XU1118 VSS VDD rst_n n899 INVx8_ASAP7_75t_R
XU1119 VSS VDD rst_n n900 INVx8_ASAP7_75t_R
XU1120 VSS VDD rst_n n901 INVx8_ASAP7_75t_R
XU1121 VSS VDD rst_n n902 INVx8_ASAP7_75t_R
XU1122 VSS VDD rst_n n903 INVx8_ASAP7_75t_R
XU1123 VSS VDD rst_n n904 INVx8_ASAP7_75t_R
XU1124 VSS VDD rst_n n905 INVx8_ASAP7_75t_R
XU1125 VSS VDD rst_n n906 INVx8_ASAP7_75t_R
XU1126 VSS VDD rst_n n907 INVx8_ASAP7_75t_R
XU1127 VSS VDD rst_n n908 INVx8_ASAP7_75t_R
XU1128 VSS VDD rst_n n909 INVx8_ASAP7_75t_R
XU1142 VSS VDD rst_n n918 INVx8_ASAP7_75t_R
XU1143 VSS VDD rst_n n919 INVx8_ASAP7_75t_R
XU1144 VSS VDD rst_n n920 INVx8_ASAP7_75t_R
XU1145 VSS VDD rst_n n921 INVx8_ASAP7_75t_R
XU1146 VSS VDD rst_n n922 INVx8_ASAP7_75t_R
XU1147 VSS VDD rst_n n923 INVx8_ASAP7_75t_R
XU1148 VSS VDD rst_n n924 INVx8_ASAP7_75t_R
XU1149 VSS VDD rst_n n925 INVx8_ASAP7_75t_R
XU1150 VSS VDD rst_n n926 INVx8_ASAP7_75t_R
XU1151 VSS VDD rst_n n927 INVx8_ASAP7_75t_R
XU1152 VSS VDD rst_n n928 INVx8_ASAP7_75t_R
XU1153 VSS VDD rst_n n929 INVx8_ASAP7_75t_R
XU1154 VSS VDD rst_n n930 INVx8_ASAP7_75t_R
XU1155 VSS VDD rst_n n931 INVx8_ASAP7_75t_R
XU1156 VSS VDD rst_n n932 INVx8_ASAP7_75t_R
XU1186 VSS VDD rst_n n937 INVx8_ASAP7_75t_R
XU1187 VSS VDD rst_n n938 INVx8_ASAP7_75t_R
XU1188 VSS VDD rst_n n939 INVx8_ASAP7_75t_R
XU1189 VSS VDD rst_n n940 INVx8_ASAP7_75t_R
XU1190 VSS VDD rst_n n941 INVx8_ASAP7_75t_R
XU1191 VSS VDD rst_n n942 INVx8_ASAP7_75t_R
XU1192 VSS VDD rst_n n943 INVx8_ASAP7_75t_R
XU1193 VSS VDD rst_n n944 INVx8_ASAP7_75t_R
XU1194 VSS VDD rst_n n945 INVx8_ASAP7_75t_R
XU1195 VSS VDD rst_n n946 INVx8_ASAP7_75t_R
XU1196 VSS VDD rst_n n947 INVx8_ASAP7_75t_R
XU1197 VSS VDD rst_n n948 INVx8_ASAP7_75t_R
XU1198 VSS VDD rst_n n949 INVx8_ASAP7_75t_R
XU1199 VSS VDD rst_n n950 INVx8_ASAP7_75t_R
XU1200 VSS VDD rst_n n951 INVx8_ASAP7_75t_R
XU1201 VSS VDD rst_n n952 INVx8_ASAP7_75t_R
XU1202 VSS VDD rst_n n953 INVx8_ASAP7_75t_R
XU1203 VSS VDD rst_n n954 INVx8_ASAP7_75t_R
XU1227 VSS VDD rst_n n958 INVx8_ASAP7_75t_R
XU1228 VSS VDD rst_n n959 INVx8_ASAP7_75t_R
XU1235 VSS VDD rst_n n962 INVx8_ASAP7_75t_R
XU1236 VSS VDD rst_n n963 INVx8_ASAP7_75t_R
XU1237 VSS VDD rst_n n972 INVx8_ASAP7_75t_R
XU1238 VSS VDD rst_n n973 INVx8_ASAP7_75t_R
XU1239 VSS VDD rst_n n976 INVx8_ASAP7_75t_R
XU1240 VSS VDD rst_n n977 INVx8_ASAP7_75t_R
XU1241 VSS VDD rst_n n978 INVx8_ASAP7_75t_R
XU1242 VSS VDD rst_n n979 INVx8_ASAP7_75t_R
XU1243 VSS VDD rst_n n980 INVx8_ASAP7_75t_R
XU1244 VSS VDD rst_n n981 INVx8_ASAP7_75t_R
XU1246 VSS VDD rst_n n982 INVx8_ASAP7_75t_R
XU1247 VSS VDD rst_n n983 INVx8_ASAP7_75t_R
XU1253 VSS VDD rst_n n985 INVx8_ASAP7_75t_R
XU1254 VSS VDD rst_n n986 INVx8_ASAP7_75t_R
XU1255 VSS VDD rst_n n987 INVx8_ASAP7_75t_R
XU1256 VSS VDD rst_n n988 INVx8_ASAP7_75t_R
XU1257 VSS VDD rst_n n1001 INVx8_ASAP7_75t_R
XU1258 VSS VDD rst_n n1006 INVx8_ASAP7_75t_R
XU1259 VSS VDD rst_n n1007 INVx8_ASAP7_75t_R
XU1260 VSS VDD rst_n n1008 INVx8_ASAP7_75t_R
XU1261 VSS VDD rst_n n1009 INVx8_ASAP7_75t_R
XU1262 VSS VDD rst_n n1010 INVx8_ASAP7_75t_R
XU1263 VSS VDD rst_n n1011 INVx8_ASAP7_75t_R
XU1264 VSS VDD rst_n n1012 INVx8_ASAP7_75t_R
XU1265 VSS VDD rst_n n1013 INVx8_ASAP7_75t_R
XU1266 VSS VDD rst_n n1014 INVx8_ASAP7_75t_R
XU1267 VSS VDD rst_n n1015 INVx8_ASAP7_75t_R
XU1268 VSS VDD rst_n n1018 INVx8_ASAP7_75t_R
XU1269 VSS VDD in_data1[127] n857 INVx8_ASAP7_75t_R
XU1270 VSS VDD in_data1[126] n856 INVx8_ASAP7_75t_R
XU1271 VSS VDD in_data1[125] n855 INVx8_ASAP7_75t_R
XU1272 VSS VDD in_data1[124] n854 INVx8_ASAP7_75t_R
XU1273 VSS VDD in_data1[123] n853 INVx8_ASAP7_75t_R
XU1274 VSS VDD in_data1[122] n852 INVx8_ASAP7_75t_R
XU1275 VSS VDD in_data1[121] n851 INVx8_ASAP7_75t_R
XU1276 VSS VDD in_data1[120] n850 INVx8_ASAP7_75t_R
XU1277 VSS VDD in_data1[119] n849 INVx8_ASAP7_75t_R
XU1278 VSS VDD in_data1[118] n848 INVx8_ASAP7_75t_R
XU1279 VSS VDD in_data1[117] n847 INVx8_ASAP7_75t_R
XU1280 VSS VDD in_data1[116] n846 INVx8_ASAP7_75t_R
XU1281 VSS VDD in_data1[115] n845 INVx8_ASAP7_75t_R
XU1282 VSS VDD in_data1[114] n844 INVx8_ASAP7_75t_R
XU1283 VSS VDD in_data1[113] n843 INVx8_ASAP7_75t_R
XU1284 VSS VDD in_data1[112] n842 INVx8_ASAP7_75t_R
XU1285 VSS VDD in_data1[111] n841 INVx8_ASAP7_75t_R
XU1286 VSS VDD in_data1[110] n840 INVx8_ASAP7_75t_R
XU1287 VSS VDD in_data1[109] n839 INVx8_ASAP7_75t_R
XU1288 VSS VDD in_data1[108] n838 INVx8_ASAP7_75t_R
XU1289 VSS VDD in_data1[107] n837 INVx8_ASAP7_75t_R
XU1290 VSS VDD in_data1[106] n836 INVx8_ASAP7_75t_R
XU1291 VSS VDD in_data1[105] n835 INVx8_ASAP7_75t_R
XU1292 VSS VDD in_data1[104] n834 INVx8_ASAP7_75t_R
XU1293 VSS VDD in_data1[103] n833 INVx8_ASAP7_75t_R
XU1294 VSS VDD in_data1[102] n832 INVx8_ASAP7_75t_R
XU1295 VSS VDD in_data1[101] n831 INVx8_ASAP7_75t_R
XU1296 VSS VDD in_data1[100] n830 INVx8_ASAP7_75t_R
XU1297 VSS VDD in_data1[99] n829 INVx8_ASAP7_75t_R
XU1298 VSS VDD in_data1[98] n828 INVx8_ASAP7_75t_R
XU1299 VSS VDD in_data1[97] n827 INVx8_ASAP7_75t_R
XU1300 VSS VDD in_data1[96] n826 INVx8_ASAP7_75t_R
XU1301 VSS VDD in_data1[95] n825 INVx8_ASAP7_75t_R
XU1302 VSS VDD in_data1[94] n824 INVx8_ASAP7_75t_R
XU1303 VSS VDD in_data1[93] n823 INVx8_ASAP7_75t_R
XU1304 VSS VDD in_data1[92] n822 INVx8_ASAP7_75t_R
XU1305 VSS VDD in_data1[91] n821 INVx8_ASAP7_75t_R
XU1306 VSS VDD in_data1[90] n820 INVx8_ASAP7_75t_R
XU1307 VSS VDD in_data1[89] n819 INVx8_ASAP7_75t_R
XU1308 VSS VDD in_data1[88] n818 INVx8_ASAP7_75t_R
XU1309 VSS VDD in_data1[87] n817 INVx8_ASAP7_75t_R
XU1310 VSS VDD in_data1[86] n816 INVx8_ASAP7_75t_R
XU1311 VSS VDD in_data1[85] n815 INVx8_ASAP7_75t_R
XU1312 VSS VDD in_data1[84] n814 INVx8_ASAP7_75t_R
XU1313 VSS VDD in_data1[83] n813 INVx8_ASAP7_75t_R
XU1314 VSS VDD in_data1[82] n812 INVx8_ASAP7_75t_R
XU1315 VSS VDD in_data1[81] n811 INVx8_ASAP7_75t_R
XU1316 VSS VDD in_data1[80] n810 INVx8_ASAP7_75t_R
XU1317 VSS VDD in_data1[79] n809 INVx8_ASAP7_75t_R
XU1318 VSS VDD in_data1[78] n808 INVx8_ASAP7_75t_R
XU1319 VSS VDD in_data1[77] n807 INVx8_ASAP7_75t_R
XU1320 VSS VDD in_data1[76] n806 INVx8_ASAP7_75t_R
XU1321 VSS VDD in_data1[75] n805 INVx8_ASAP7_75t_R
XU1322 VSS VDD in_data1[74] n804 INVx8_ASAP7_75t_R
XU1323 VSS VDD in_data1[73] n803 INVx8_ASAP7_75t_R
XU1324 VSS VDD in_data1[72] n802 INVx8_ASAP7_75t_R
XU1325 VSS VDD in_data1[71] n801 INVx8_ASAP7_75t_R
XU1326 VSS VDD in_data1[70] n800 INVx8_ASAP7_75t_R
XU1327 VSS VDD in_data1[69] n799 INVx8_ASAP7_75t_R
XU1328 VSS VDD in_data1[68] n798 INVx8_ASAP7_75t_R
XU1329 VSS VDD in_data1[67] n797 INVx8_ASAP7_75t_R
XU1330 VSS VDD in_data1[66] n796 INVx8_ASAP7_75t_R
XU1331 VSS VDD in_data1[65] n795 INVx8_ASAP7_75t_R
XU1332 VSS VDD in_data1[64] n794 INVx8_ASAP7_75t_R
XU1333 VSS VDD in_data1[63] n793 INVx8_ASAP7_75t_R
XU1334 VSS VDD in_data1[62] n792 INVx8_ASAP7_75t_R
XU1335 VSS VDD in_data1[61] n791 INVx8_ASAP7_75t_R
XU1336 VSS VDD in_data1[60] n790 INVx8_ASAP7_75t_R
XU1337 VSS VDD in_data1[59] n789 INVx8_ASAP7_75t_R
XU1338 VSS VDD in_data1[58] n788 INVx8_ASAP7_75t_R
XU1339 VSS VDD in_data1[57] n787 INVx8_ASAP7_75t_R
XU1340 VSS VDD in_data1[56] n786 INVx8_ASAP7_75t_R
XU1341 VSS VDD in_data1[55] n785 INVx8_ASAP7_75t_R
XU1342 VSS VDD in_data1[54] n784 INVx8_ASAP7_75t_R
XU1343 VSS VDD in_data1[53] n783 INVx8_ASAP7_75t_R
XU1344 VSS VDD in_data1[52] n782 INVx8_ASAP7_75t_R
XU1345 VSS VDD in_data1[51] n781 INVx8_ASAP7_75t_R
XU1346 VSS VDD in_data1[50] n780 INVx8_ASAP7_75t_R
XU1347 VSS VDD in_data1[49] n779 INVx8_ASAP7_75t_R
XU1348 VSS VDD in_data1[48] n778 INVx8_ASAP7_75t_R
XU1349 VSS VDD in_data1[47] n777 INVx8_ASAP7_75t_R
XU1350 VSS VDD in_data1[46] n776 INVx8_ASAP7_75t_R
XU1351 VSS VDD in_data1[45] n775 INVx8_ASAP7_75t_R
XU1352 VSS VDD in_data1[44] n774 INVx8_ASAP7_75t_R
XU1353 VSS VDD in_data1[43] n773 INVx8_ASAP7_75t_R
XU1354 VSS VDD in_data1[42] n772 INVx8_ASAP7_75t_R
XU1355 VSS VDD in_data1[41] n771 INVx8_ASAP7_75t_R
XU1356 VSS VDD in_data1[40] n770 INVx8_ASAP7_75t_R
XU1357 VSS VDD in_data1[39] n769 INVx8_ASAP7_75t_R
XU1358 VSS VDD in_data1[38] n768 INVx8_ASAP7_75t_R
XU1359 VSS VDD in_data1[37] n767 INVx8_ASAP7_75t_R
XU1360 VSS VDD in_data1[36] n766 INVx8_ASAP7_75t_R
XU1361 VSS VDD in_data1[35] n765 INVx8_ASAP7_75t_R
XU1362 VSS VDD in_data1[34] n764 INVx8_ASAP7_75t_R
XU1363 VSS VDD in_data1[33] n763 INVx8_ASAP7_75t_R
XU1364 VSS VDD in_data1[32] n762 INVx8_ASAP7_75t_R
XU1365 VSS VDD in_data1[31] n761 INVx8_ASAP7_75t_R
XU1366 VSS VDD in_data1[30] n760 INVx8_ASAP7_75t_R
XU1367 VSS VDD in_data1[29] n759 INVx8_ASAP7_75t_R
XU1368 VSS VDD in_data1[28] n758 INVx8_ASAP7_75t_R
XU1369 VSS VDD in_data1[27] n757 INVx8_ASAP7_75t_R
XU1370 VSS VDD in_data1[26] n756 INVx8_ASAP7_75t_R
XU1371 VSS VDD in_data1[25] n755 INVx8_ASAP7_75t_R
XU1372 VSS VDD in_data1[24] n754 INVx8_ASAP7_75t_R
XU1373 VSS VDD in_data1[23] n753 INVx8_ASAP7_75t_R
XU1374 VSS VDD in_data1[22] n752 INVx8_ASAP7_75t_R
XU1375 VSS VDD in_data1[21] n751 INVx8_ASAP7_75t_R
XU1376 VSS VDD in_data1[20] n750 INVx8_ASAP7_75t_R
XU1377 VSS VDD in_data1[19] n749 INVx8_ASAP7_75t_R
XU1378 VSS VDD in_data1[18] n748 INVx8_ASAP7_75t_R
XU1379 VSS VDD in_data1[17] n747 INVx8_ASAP7_75t_R
XU1380 VSS VDD in_data1[16] n746 INVx8_ASAP7_75t_R
XU1381 VSS VDD in_data1[15] n745 INVx8_ASAP7_75t_R
XU1382 VSS VDD in_data1[14] n744 INVx8_ASAP7_75t_R
XU1383 VSS VDD in_data1[13] n743 INVx8_ASAP7_75t_R
XU1384 VSS VDD in_data1[12] n742 INVx8_ASAP7_75t_R
XU1385 VSS VDD in_data1[11] n741 INVx8_ASAP7_75t_R
XU1386 VSS VDD in_data1[10] n740 INVx8_ASAP7_75t_R
XU1387 VSS VDD in_data1[9] n739 INVx8_ASAP7_75t_R
XU1388 VSS VDD in_data1[8] n738 INVx8_ASAP7_75t_R
XU1389 VSS VDD in_data1[7] n737 INVx8_ASAP7_75t_R
XU1390 VSS VDD in_data1[6] n736 INVx8_ASAP7_75t_R
XU1391 VSS VDD in_data1[5] n735 INVx8_ASAP7_75t_R
XU1392 VSS VDD in_data1[4] n734 INVx8_ASAP7_75t_R
XU1393 VSS VDD in_data1[3] n733 INVx8_ASAP7_75t_R
XU1394 VSS VDD in_data1[2] n732 INVx8_ASAP7_75t_R
XU1395 VSS VDD in_data1[1] n731 INVx8_ASAP7_75t_R
XU1396 VSS VDD in_data1[0] n730 INVx8_ASAP7_75t_R
XU1397 VSS VDD in_data2[127] n729 INVx8_ASAP7_75t_R
XU1398 VSS VDD in_data2[126] n728 INVx8_ASAP7_75t_R
XU1399 VSS VDD in_data2[125] n727 INVx8_ASAP7_75t_R
XU1400 VSS VDD in_data2[124] n726 INVx8_ASAP7_75t_R
XU1401 VSS VDD in_data2[123] n725 INVx8_ASAP7_75t_R
XU1402 VSS VDD in_data2[122] n724 INVx8_ASAP7_75t_R
XU1403 VSS VDD in_data2[121] n723 INVx8_ASAP7_75t_R
XU1404 VSS VDD in_data2[120] n722 INVx8_ASAP7_75t_R
XU1405 VSS VDD in_data2[119] n721 INVx8_ASAP7_75t_R
XU1406 VSS VDD in_data2[118] n720 INVx8_ASAP7_75t_R
XU1407 VSS VDD in_data2[117] n719 INVx8_ASAP7_75t_R
XU1408 VSS VDD in_data2[116] n718 INVx8_ASAP7_75t_R
XU1409 VSS VDD in_data2[115] n717 INVx8_ASAP7_75t_R
XU1410 VSS VDD in_data2[114] n716 INVx8_ASAP7_75t_R
XU1411 VSS VDD in_data2[113] n715 INVx8_ASAP7_75t_R
XU1412 VSS VDD in_data2[112] n714 INVx8_ASAP7_75t_R
XU1413 VSS VDD in_data2[111] n713 INVx8_ASAP7_75t_R
XU1414 VSS VDD in_data2[110] n712 INVx8_ASAP7_75t_R
XU1415 VSS VDD in_data2[109] n711 INVx8_ASAP7_75t_R
XU1416 VSS VDD in_data2[108] n710 INVx8_ASAP7_75t_R
XU1417 VSS VDD in_data2[107] n709 INVx8_ASAP7_75t_R
XU1418 VSS VDD in_data2[106] n708 INVx8_ASAP7_75t_R
XU1419 VSS VDD in_data2[105] n707 INVx8_ASAP7_75t_R
XU1420 VSS VDD in_data2[104] n706 INVx8_ASAP7_75t_R
XU1421 VSS VDD in_data2[103] n705 INVx8_ASAP7_75t_R
XU1422 VSS VDD in_data2[102] n704 INVx8_ASAP7_75t_R
XU1423 VSS VDD in_data2[101] n703 INVx8_ASAP7_75t_R
XU1424 VSS VDD in_data2[100] n702 INVx8_ASAP7_75t_R
XU1425 VSS VDD in_data2[99] n701 INVx8_ASAP7_75t_R
XU1426 VSS VDD in_data2[98] n700 INVx8_ASAP7_75t_R
XU1427 VSS VDD in_data2[97] n699 INVx8_ASAP7_75t_R
XU1428 VSS VDD in_data2[96] n698 INVx8_ASAP7_75t_R
XU1429 VSS VDD in_data2[95] n697 INVx8_ASAP7_75t_R
XU1430 VSS VDD in_data2[94] n696 INVx8_ASAP7_75t_R
XU1431 VSS VDD in_data2[93] n695 INVx8_ASAP7_75t_R
XU1432 VSS VDD in_data2[92] n694 INVx8_ASAP7_75t_R
XU1433 VSS VDD in_data2[91] n693 INVx8_ASAP7_75t_R
XU1434 VSS VDD in_data2[90] n692 INVx8_ASAP7_75t_R
XU1435 VSS VDD in_data2[89] n691 INVx8_ASAP7_75t_R
XU1436 VSS VDD in_data2[88] n690 INVx8_ASAP7_75t_R
XU1437 VSS VDD in_data2[87] n689 INVx8_ASAP7_75t_R
XU1438 VSS VDD in_data2[86] n688 INVx8_ASAP7_75t_R
XU1439 VSS VDD in_data2[85] n687 INVx8_ASAP7_75t_R
XU1440 VSS VDD in_data2[84] n686 INVx8_ASAP7_75t_R
XU1441 VSS VDD in_data2[83] n685 INVx8_ASAP7_75t_R
XU1442 VSS VDD in_data2[82] n684 INVx8_ASAP7_75t_R
XU1443 VSS VDD in_data2[81] n683 INVx8_ASAP7_75t_R
XU1444 VSS VDD in_data2[80] n682 INVx8_ASAP7_75t_R
XU1445 VSS VDD in_data2[79] n681 INVx8_ASAP7_75t_R
XU1446 VSS VDD in_data2[78] n680 INVx8_ASAP7_75t_R
XU1447 VSS VDD in_data2[77] n679 INVx8_ASAP7_75t_R
XU1448 VSS VDD in_data2[76] n678 INVx8_ASAP7_75t_R
XU1449 VSS VDD in_data2[75] n677 INVx8_ASAP7_75t_R
XU1450 VSS VDD in_data2[74] n676 INVx8_ASAP7_75t_R
XU1451 VSS VDD in_data2[73] n675 INVx8_ASAP7_75t_R
XU1452 VSS VDD in_data2[72] n674 INVx8_ASAP7_75t_R
XU1453 VSS VDD in_data2[71] n673 INVx8_ASAP7_75t_R
XU1454 VSS VDD in_data2[70] n672 INVx8_ASAP7_75t_R
XU1455 VSS VDD in_data2[69] n671 INVx8_ASAP7_75t_R
XU1456 VSS VDD in_data2[68] n670 INVx8_ASAP7_75t_R
XU1457 VSS VDD in_data2[67] n669 INVx8_ASAP7_75t_R
XU1458 VSS VDD in_data2[66] n668 INVx8_ASAP7_75t_R
XU1459 VSS VDD in_data2[65] n667 INVx8_ASAP7_75t_R
XU1460 VSS VDD in_data2[64] n666 INVx8_ASAP7_75t_R
XU1461 VSS VDD in_data2[63] n665 INVx8_ASAP7_75t_R
XU1462 VSS VDD in_data2[62] n664 INVx8_ASAP7_75t_R
XU1463 VSS VDD in_data2[61] n663 INVx8_ASAP7_75t_R
XU1464 VSS VDD in_data2[60] n662 INVx8_ASAP7_75t_R
XU1465 VSS VDD in_data2[59] n661 INVx8_ASAP7_75t_R
XU1466 VSS VDD in_data2[58] n660 INVx8_ASAP7_75t_R
XU1467 VSS VDD in_data2[57] n659 INVx8_ASAP7_75t_R
XU1468 VSS VDD in_data2[56] n658 INVx8_ASAP7_75t_R
XU1469 VSS VDD in_data2[55] n657 INVx8_ASAP7_75t_R
XU1470 VSS VDD in_data2[54] n656 INVx8_ASAP7_75t_R
XU1471 VSS VDD in_data2[53] n655 INVx8_ASAP7_75t_R
XU1472 VSS VDD in_data2[52] n654 INVx8_ASAP7_75t_R
XU1473 VSS VDD in_data2[51] n653 INVx8_ASAP7_75t_R
XU1474 VSS VDD in_data2[50] n652 INVx8_ASAP7_75t_R
XU1475 VSS VDD in_data2[49] n651 INVx8_ASAP7_75t_R
XU1476 VSS VDD in_data2[48] n650 INVx8_ASAP7_75t_R
XU1477 VSS VDD in_data2[47] n649 INVx8_ASAP7_75t_R
XU1478 VSS VDD in_data2[46] n648 INVx8_ASAP7_75t_R
XU1479 VSS VDD in_data2[45] n647 INVx8_ASAP7_75t_R
XU1480 VSS VDD in_data2[44] n646 INVx8_ASAP7_75t_R
XU1481 VSS VDD in_data2[43] n645 INVx8_ASAP7_75t_R
XU1482 VSS VDD in_data2[42] n644 INVx8_ASAP7_75t_R
XU1483 VSS VDD in_data2[41] n643 INVx8_ASAP7_75t_R
XU1484 VSS VDD in_data2[40] n642 INVx8_ASAP7_75t_R
XU1485 VSS VDD in_data2[39] n641 INVx8_ASAP7_75t_R
XU1486 VSS VDD in_data2[38] n640 INVx8_ASAP7_75t_R
XU1487 VSS VDD in_data2[37] n639 INVx8_ASAP7_75t_R
XU1488 VSS VDD in_data2[36] n638 INVx8_ASAP7_75t_R
XU1489 VSS VDD in_data2[35] n637 INVx8_ASAP7_75t_R
XU1490 VSS VDD in_data2[34] n636 INVx8_ASAP7_75t_R
XU1491 VSS VDD in_data2[33] n635 INVx8_ASAP7_75t_R
XU1492 VSS VDD in_data2[32] n634 INVx8_ASAP7_75t_R
XU1493 VSS VDD in_data2[31] n633 INVx8_ASAP7_75t_R
XU1494 VSS VDD in_data2[30] n632 INVx8_ASAP7_75t_R
XU1495 VSS VDD in_data2[29] n631 INVx8_ASAP7_75t_R
XU1496 VSS VDD in_data2[28] n630 INVx8_ASAP7_75t_R
XU1497 VSS VDD in_data2[27] n629 INVx8_ASAP7_75t_R
XU1498 VSS VDD in_data2[26] n628 INVx8_ASAP7_75t_R
XU1499 VSS VDD in_data2[25] n627 INVx8_ASAP7_75t_R
XU1500 VSS VDD in_data2[24] n626 INVx8_ASAP7_75t_R
XU1501 VSS VDD in_data2[23] n625 INVx8_ASAP7_75t_R
XU1502 VSS VDD in_data2[22] n624 INVx8_ASAP7_75t_R
XU1503 VSS VDD in_data2[21] n623 INVx8_ASAP7_75t_R
XU1504 VSS VDD in_data2[20] n622 INVx8_ASAP7_75t_R
XU1505 VSS VDD in_data2[19] n621 INVx8_ASAP7_75t_R
XU1506 VSS VDD in_data2[18] n620 INVx8_ASAP7_75t_R
XU1507 VSS VDD in_data2[17] n619 INVx8_ASAP7_75t_R
XU1508 VSS VDD in_data2[16] n618 INVx8_ASAP7_75t_R
XU1509 VSS VDD in_data2[15] n617 INVx8_ASAP7_75t_R
XU1510 VSS VDD in_data2[14] n616 INVx8_ASAP7_75t_R
XU1511 VSS VDD in_data2[13] n615 INVx8_ASAP7_75t_R
XU1512 VSS VDD in_data2[12] n614 INVx8_ASAP7_75t_R
XU1513 VSS VDD in_data2[11] n613 INVx8_ASAP7_75t_R
XU1514 VSS VDD in_data2[10] n612 INVx8_ASAP7_75t_R
XU1515 VSS VDD in_data2[9] n611 INVx8_ASAP7_75t_R
XU1516 VSS VDD in_data2[8] n610 INVx8_ASAP7_75t_R
XU1517 VSS VDD in_data2[7] n609 INVx8_ASAP7_75t_R
XU1518 VSS VDD in_data2[6] n608 INVx8_ASAP7_75t_R
XU1519 VSS VDD in_data2[5] n607 INVx8_ASAP7_75t_R
XU1520 VSS VDD in_data2[4] n606 INVx8_ASAP7_75t_R
XU1521 VSS VDD in_data2[3] n605 INVx8_ASAP7_75t_R
XU1522 VSS VDD in_data2[2] n604 INVx8_ASAP7_75t_R
XU1523 VSS VDD in_data2[1] n603 INVx8_ASAP7_75t_R
XU1524 VSS VDD in_data2[0] n602 INVx8_ASAP7_75t_R
XU1525 VSS VDD in_data3[127] n601 INVx8_ASAP7_75t_R
XU1526 VSS VDD in_data3[126] n600 INVx8_ASAP7_75t_R
XU1527 VSS VDD in_data3[125] n599 INVx8_ASAP7_75t_R
XU1528 VSS VDD in_data3[124] n598 INVx8_ASAP7_75t_R
XU1529 VSS VDD in_data3[123] n597 INVx8_ASAP7_75t_R
XU1530 VSS VDD in_data3[122] n596 INVx8_ASAP7_75t_R
XU1531 VSS VDD in_data3[121] n595 INVx8_ASAP7_75t_R
XU1532 VSS VDD in_data3[120] n594 INVx8_ASAP7_75t_R
XU1533 VSS VDD in_data3[119] n593 INVx8_ASAP7_75t_R
XU1534 VSS VDD in_data3[118] n592 INVx8_ASAP7_75t_R
XU1535 VSS VDD in_data3[117] n591 INVx8_ASAP7_75t_R
XU1536 VSS VDD in_data3[116] n590 INVx8_ASAP7_75t_R
XU1537 VSS VDD in_data3[115] n589 INVx8_ASAP7_75t_R
XU1538 VSS VDD in_data3[114] n588 INVx8_ASAP7_75t_R
XU1539 VSS VDD in_data3[113] n587 INVx8_ASAP7_75t_R
XU1540 VSS VDD in_data3[112] n586 INVx8_ASAP7_75t_R
XU1541 VSS VDD in_data3[111] n585 INVx8_ASAP7_75t_R
XU1542 VSS VDD in_data3[110] n584 INVx8_ASAP7_75t_R
XU1543 VSS VDD in_data3[109] n583 INVx8_ASAP7_75t_R
XU1544 VSS VDD in_data3[108] n582 INVx8_ASAP7_75t_R
XU1545 VSS VDD in_data3[107] n581 INVx8_ASAP7_75t_R
XU1546 VSS VDD in_data3[106] n580 INVx8_ASAP7_75t_R
XU1547 VSS VDD in_data3[105] n579 INVx8_ASAP7_75t_R
XU1548 VSS VDD in_data3[104] n578 INVx8_ASAP7_75t_R
XU1549 VSS VDD in_data3[103] n577 INVx8_ASAP7_75t_R
XU1550 VSS VDD in_data3[102] n576 INVx8_ASAP7_75t_R
XU1551 VSS VDD in_data3[101] n575 INVx8_ASAP7_75t_R
XU1552 VSS VDD in_data3[100] n574 INVx8_ASAP7_75t_R
XU1553 VSS VDD in_data3[99] n573 INVx8_ASAP7_75t_R
XU1554 VSS VDD in_data3[98] n572 INVx8_ASAP7_75t_R
XU1555 VSS VDD in_data3[97] n571 INVx8_ASAP7_75t_R
XU1556 VSS VDD in_data3[96] n570 INVx8_ASAP7_75t_R
XU1557 VSS VDD in_data3[95] n569 INVx8_ASAP7_75t_R
XU1558 VSS VDD in_data3[94] n568 INVx8_ASAP7_75t_R
XU1559 VSS VDD in_data3[93] n567 INVx8_ASAP7_75t_R
XU1560 VSS VDD in_data3[92] n566 INVx8_ASAP7_75t_R
XU1561 VSS VDD in_data3[91] n565 INVx8_ASAP7_75t_R
XU1562 VSS VDD in_data3[90] n564 INVx8_ASAP7_75t_R
XU1563 VSS VDD in_data3[89] n563 INVx8_ASAP7_75t_R
XU1564 VSS VDD in_data3[88] n562 INVx8_ASAP7_75t_R
XU1565 VSS VDD in_data3[87] n561 INVx8_ASAP7_75t_R
XU1566 VSS VDD in_data3[86] n560 INVx8_ASAP7_75t_R
XU1567 VSS VDD in_data3[85] n559 INVx8_ASAP7_75t_R
XU1568 VSS VDD in_data3[84] n558 INVx8_ASAP7_75t_R
XU1569 VSS VDD in_data3[83] n557 INVx8_ASAP7_75t_R
XU1570 VSS VDD in_data3[82] n556 INVx8_ASAP7_75t_R
XU1571 VSS VDD in_data3[81] n555 INVx8_ASAP7_75t_R
XU1572 VSS VDD in_data3[80] n554 INVx8_ASAP7_75t_R
XU1573 VSS VDD in_data3[79] n553 INVx8_ASAP7_75t_R
XU1574 VSS VDD in_data3[78] n552 INVx8_ASAP7_75t_R
XU1575 VSS VDD in_data3[77] n551 INVx8_ASAP7_75t_R
XU1576 VSS VDD in_data3[76] n550 INVx8_ASAP7_75t_R
XU1577 VSS VDD in_data3[75] n549 INVx8_ASAP7_75t_R
XU1578 VSS VDD in_data3[74] n548 INVx8_ASAP7_75t_R
XU1579 VSS VDD in_data3[73] n547 INVx8_ASAP7_75t_R
XU1580 VSS VDD in_data3[72] n546 INVx8_ASAP7_75t_R
XU1581 VSS VDD in_data3[71] n545 INVx8_ASAP7_75t_R
XU1582 VSS VDD in_data3[70] n544 INVx8_ASAP7_75t_R
XU1583 VSS VDD in_data3[69] n543 INVx8_ASAP7_75t_R
XU1584 VSS VDD in_data3[68] n542 INVx8_ASAP7_75t_R
XU1585 VSS VDD in_data3[67] n541 INVx8_ASAP7_75t_R
XU1586 VSS VDD in_data3[66] n540 INVx8_ASAP7_75t_R
XU1587 VSS VDD in_data3[65] n539 INVx8_ASAP7_75t_R
XU1588 VSS VDD in_data3[64] n538 INVx8_ASAP7_75t_R
XU1589 VSS VDD in_data3[63] n537 INVx8_ASAP7_75t_R
XU1590 VSS VDD in_data3[62] n536 INVx8_ASAP7_75t_R
XU1591 VSS VDD in_data3[61] n535 INVx8_ASAP7_75t_R
XU1592 VSS VDD in_data3[60] n534 INVx8_ASAP7_75t_R
XU1593 VSS VDD in_data3[59] n533 INVx8_ASAP7_75t_R
XU1594 VSS VDD in_data3[58] n532 INVx8_ASAP7_75t_R
XU1595 VSS VDD in_data3[57] n531 INVx8_ASAP7_75t_R
XU1596 VSS VDD in_data3[56] n530 INVx8_ASAP7_75t_R
XU1597 VSS VDD in_data3[55] n529 INVx8_ASAP7_75t_R
XU1598 VSS VDD in_data3[54] n528 INVx8_ASAP7_75t_R
XU1599 VSS VDD in_data3[53] n527 INVx8_ASAP7_75t_R
XU1600 VSS VDD in_data3[52] n526 INVx8_ASAP7_75t_R
XU1601 VSS VDD in_data3[51] n525 INVx8_ASAP7_75t_R
XU1602 VSS VDD in_data3[50] n524 INVx8_ASAP7_75t_R
XU1603 VSS VDD in_data3[49] n523 INVx8_ASAP7_75t_R
XU1604 VSS VDD in_data3[48] n522 INVx8_ASAP7_75t_R
XU1605 VSS VDD in_data3[47] n521 INVx8_ASAP7_75t_R
XU1606 VSS VDD in_data3[46] n520 INVx8_ASAP7_75t_R
XU1607 VSS VDD in_data3[45] n519 INVx8_ASAP7_75t_R
XU1608 VSS VDD in_data3[44] n518 INVx8_ASAP7_75t_R
XU1609 VSS VDD in_data3[43] n517 INVx8_ASAP7_75t_R
XU1610 VSS VDD in_data3[42] n516 INVx8_ASAP7_75t_R
XU1611 VSS VDD in_data3[41] n515 INVx8_ASAP7_75t_R
XU1612 VSS VDD in_data3[40] n514 INVx8_ASAP7_75t_R
XU1613 VSS VDD in_data3[39] n513 INVx8_ASAP7_75t_R
XU1614 VSS VDD in_data3[38] n512 INVx8_ASAP7_75t_R
XU1615 VSS VDD in_data3[37] n511 INVx8_ASAP7_75t_R
XU1616 VSS VDD in_data3[36] n510 INVx8_ASAP7_75t_R
XU1617 VSS VDD in_data3[35] n509 INVx8_ASAP7_75t_R
XU1618 VSS VDD in_data3[34] n508 INVx8_ASAP7_75t_R
XU1619 VSS VDD in_data3[33] n507 INVx8_ASAP7_75t_R
XU1620 VSS VDD in_data3[32] n506 INVx8_ASAP7_75t_R
XU1621 VSS VDD in_data3[31] n505 INVx8_ASAP7_75t_R
XU1622 VSS VDD in_data3[30] n504 INVx8_ASAP7_75t_R
XU1623 VSS VDD in_data3[29] n503 INVx8_ASAP7_75t_R
XU1624 VSS VDD in_data3[28] n502 INVx8_ASAP7_75t_R
XU1625 VSS VDD in_data3[27] n501 INVx8_ASAP7_75t_R
XU1626 VSS VDD in_data3[26] n500 INVx8_ASAP7_75t_R
XU1627 VSS VDD in_data3[25] n499 INVx8_ASAP7_75t_R
XU1628 VSS VDD in_data3[24] n498 INVx8_ASAP7_75t_R
XU1629 VSS VDD in_data3[23] n497 INVx8_ASAP7_75t_R
XU1630 VSS VDD in_data3[22] n496 INVx8_ASAP7_75t_R
XU1631 VSS VDD in_data3[21] n495 INVx8_ASAP7_75t_R
XU1632 VSS VDD in_data3[20] n494 INVx8_ASAP7_75t_R
XU1633 VSS VDD in_data3[19] n493 INVx8_ASAP7_75t_R
XU1634 VSS VDD in_data3[18] n492 INVx8_ASAP7_75t_R
XU1635 VSS VDD in_data3[17] n491 INVx8_ASAP7_75t_R
XU1636 VSS VDD in_data3[16] n490 INVx8_ASAP7_75t_R
XU1637 VSS VDD in_data3[15] n489 INVx8_ASAP7_75t_R
XU1638 VSS VDD in_data3[14] n488 INVx8_ASAP7_75t_R
XU1639 VSS VDD in_data3[13] n487 INVx8_ASAP7_75t_R
XU1640 VSS VDD in_data3[12] n486 INVx8_ASAP7_75t_R
XU1641 VSS VDD in_data3[11] n485 INVx8_ASAP7_75t_R
XU1642 VSS VDD in_data3[10] n484 INVx8_ASAP7_75t_R
XU1643 VSS VDD in_data3[9] n483 INVx8_ASAP7_75t_R
XU1644 VSS VDD in_data3[8] n482 INVx8_ASAP7_75t_R
XU1645 VSS VDD in_data3[7] n481 INVx8_ASAP7_75t_R
XU1646 VSS VDD in_data3[6] n480 INVx8_ASAP7_75t_R
XU1647 VSS VDD in_data3[5] n479 INVx8_ASAP7_75t_R
XU1648 VSS VDD in_data3[4] n478 INVx8_ASAP7_75t_R
XU1649 VSS VDD in_data3[3] n477 INVx8_ASAP7_75t_R
XU1650 VSS VDD in_data3[2] n476 INVx8_ASAP7_75t_R
XU1651 VSS VDD in_data3[1] n475 INVx8_ASAP7_75t_R
XU1652 VSS VDD in_data3[0] n474 INVx8_ASAP7_75t_R
XU1653 VSS VDD in_data4[127] n473 INVx8_ASAP7_75t_R
XU1654 VSS VDD in_data4[126] n472 INVx8_ASAP7_75t_R
XU1655 VSS VDD in_data4[125] n471 INVx8_ASAP7_75t_R
XU1656 VSS VDD in_data4[124] n470 INVx8_ASAP7_75t_R
XU1657 VSS VDD in_data4[123] n469 INVx8_ASAP7_75t_R
XU1658 VSS VDD in_data4[122] n468 INVx8_ASAP7_75t_R
XU1659 VSS VDD in_data4[121] n467 INVx8_ASAP7_75t_R
XU1660 VSS VDD in_data4[120] n466 INVx8_ASAP7_75t_R
XU1661 VSS VDD in_data4[119] n465 INVx8_ASAP7_75t_R
XU1662 VSS VDD in_data4[118] n464 INVx8_ASAP7_75t_R
XU1663 VSS VDD in_data4[117] n463 INVx8_ASAP7_75t_R
XU1664 VSS VDD in_data4[116] n462 INVx8_ASAP7_75t_R
XU1665 VSS VDD in_data4[115] n461 INVx8_ASAP7_75t_R
XU1666 VSS VDD in_data4[114] n460 INVx8_ASAP7_75t_R
XU1667 VSS VDD in_data4[113] n459 INVx8_ASAP7_75t_R
XU1668 VSS VDD in_data4[112] n458 INVx8_ASAP7_75t_R
XU1669 VSS VDD in_data4[111] n457 INVx8_ASAP7_75t_R
XU1670 VSS VDD in_data4[110] n456 INVx8_ASAP7_75t_R
XU1671 VSS VDD in_data4[109] n455 INVx8_ASAP7_75t_R
XU1672 VSS VDD in_data4[108] n454 INVx8_ASAP7_75t_R
XU1673 VSS VDD in_data4[107] n453 INVx8_ASAP7_75t_R
XU1674 VSS VDD in_data4[106] n452 INVx8_ASAP7_75t_R
XU1675 VSS VDD in_data4[105] n451 INVx8_ASAP7_75t_R
XU1676 VSS VDD in_data4[104] n450 INVx8_ASAP7_75t_R
XU1677 VSS VDD in_data4[103] n449 INVx8_ASAP7_75t_R
XU1678 VSS VDD in_data4[102] n448 INVx8_ASAP7_75t_R
XU1679 VSS VDD in_data4[101] n447 INVx8_ASAP7_75t_R
XU1680 VSS VDD in_data4[100] n446 INVx8_ASAP7_75t_R
XU1681 VSS VDD in_data4[99] n445 INVx8_ASAP7_75t_R
XU1682 VSS VDD in_data4[98] n444 INVx8_ASAP7_75t_R
XU1683 VSS VDD in_data4[97] n443 INVx8_ASAP7_75t_R
XU1684 VSS VDD in_data4[96] n442 INVx8_ASAP7_75t_R
XU1685 VSS VDD in_data4[95] n441 INVx8_ASAP7_75t_R
XU1686 VSS VDD in_data4[94] n440 INVx8_ASAP7_75t_R
XU1687 VSS VDD in_data4[93] n439 INVx8_ASAP7_75t_R
XU1688 VSS VDD in_data4[92] n438 INVx8_ASAP7_75t_R
XU1689 VSS VDD in_data4[91] n437 INVx8_ASAP7_75t_R
XU1690 VSS VDD in_data4[90] n436 INVx8_ASAP7_75t_R
XU1691 VSS VDD in_data4[89] n435 INVx8_ASAP7_75t_R
XU1692 VSS VDD in_data4[88] n434 INVx8_ASAP7_75t_R
XU1693 VSS VDD in_data4[87] n433 INVx8_ASAP7_75t_R
XU1694 VSS VDD in_data4[86] n432 INVx8_ASAP7_75t_R
XU1695 VSS VDD in_data4[85] n431 INVx8_ASAP7_75t_R
XU1696 VSS VDD in_data4[84] n430 INVx8_ASAP7_75t_R
XU1697 VSS VDD in_data4[83] n429 INVx8_ASAP7_75t_R
XU1698 VSS VDD in_data4[82] n428 INVx8_ASAP7_75t_R
XU1699 VSS VDD in_data4[81] n427 INVx8_ASAP7_75t_R
XU1700 VSS VDD in_data4[80] n426 INVx8_ASAP7_75t_R
XU1701 VSS VDD in_data4[79] n425 INVx8_ASAP7_75t_R
XU1702 VSS VDD in_data4[78] n424 INVx8_ASAP7_75t_R
XU1703 VSS VDD in_data4[77] n423 INVx8_ASAP7_75t_R
XU1704 VSS VDD in_data4[76] n422 INVx8_ASAP7_75t_R
XU1705 VSS VDD in_data4[75] n421 INVx8_ASAP7_75t_R
XU1706 VSS VDD in_data4[74] n420 INVx8_ASAP7_75t_R
XU1707 VSS VDD in_data4[73] n419 INVx8_ASAP7_75t_R
XU1708 VSS VDD in_data4[72] n418 INVx8_ASAP7_75t_R
XU1709 VSS VDD in_data4[71] n417 INVx8_ASAP7_75t_R
XU1710 VSS VDD in_data4[70] n416 INVx8_ASAP7_75t_R
XU1711 VSS VDD in_data4[69] n415 INVx8_ASAP7_75t_R
XU1712 VSS VDD in_data4[68] n414 INVx8_ASAP7_75t_R
XU1713 VSS VDD in_data4[67] n413 INVx8_ASAP7_75t_R
XU1714 VSS VDD in_data4[66] n412 INVx8_ASAP7_75t_R
XU1715 VSS VDD in_data4[65] n411 INVx8_ASAP7_75t_R
XU1716 VSS VDD in_data4[64] n410 INVx8_ASAP7_75t_R
XU1717 VSS VDD in_data4[63] n409 INVx8_ASAP7_75t_R
XU1718 VSS VDD in_data4[62] n408 INVx8_ASAP7_75t_R
XU1719 VSS VDD in_data4[61] n407 INVx8_ASAP7_75t_R
XU1720 VSS VDD in_data4[60] n406 INVx8_ASAP7_75t_R
XU1721 VSS VDD in_data4[59] n405 INVx8_ASAP7_75t_R
XU1722 VSS VDD in_data4[58] n404 INVx8_ASAP7_75t_R
XU1723 VSS VDD in_data4[57] n403 INVx8_ASAP7_75t_R
XU1724 VSS VDD in_data4[56] n402 INVx8_ASAP7_75t_R
XU1725 VSS VDD in_data4[55] n401 INVx8_ASAP7_75t_R
XU1726 VSS VDD in_data4[54] n400 INVx8_ASAP7_75t_R
XU1727 VSS VDD in_data4[53] n399 INVx8_ASAP7_75t_R
XU1728 VSS VDD in_data4[52] n398 INVx8_ASAP7_75t_R
XU1729 VSS VDD in_data4[51] n397 INVx8_ASAP7_75t_R
XU1730 VSS VDD in_data4[50] n396 INVx8_ASAP7_75t_R
XU1731 VSS VDD in_data4[49] n395 INVx8_ASAP7_75t_R
XU1732 VSS VDD in_data4[48] n394 INVx8_ASAP7_75t_R
XU1733 VSS VDD in_data4[47] n393 INVx8_ASAP7_75t_R
XU1734 VSS VDD in_data4[46] n392 INVx8_ASAP7_75t_R
XU1735 VSS VDD in_data4[45] n391 INVx8_ASAP7_75t_R
XU1736 VSS VDD in_data4[44] n390 INVx8_ASAP7_75t_R
XU1737 VSS VDD in_data4[43] n389 INVx8_ASAP7_75t_R
XU1738 VSS VDD in_data4[42] n388 INVx8_ASAP7_75t_R
XU1739 VSS VDD in_data4[41] n387 INVx8_ASAP7_75t_R
XU1740 VSS VDD in_data4[40] n386 INVx8_ASAP7_75t_R
XU1741 VSS VDD in_data4[39] n385 INVx8_ASAP7_75t_R
XU1742 VSS VDD in_data4[38] n384 INVx8_ASAP7_75t_R
XU1743 VSS VDD in_data4[37] n383 INVx8_ASAP7_75t_R
XU1744 VSS VDD in_data4[36] n382 INVx8_ASAP7_75t_R
XU1745 VSS VDD in_data4[35] n381 INVx8_ASAP7_75t_R
XU1746 VSS VDD in_data4[34] n380 INVx8_ASAP7_75t_R
XU1747 VSS VDD in_data4[33] n379 INVx8_ASAP7_75t_R
XU1748 VSS VDD in_data4[32] n378 INVx8_ASAP7_75t_R
XU1749 VSS VDD in_data4[31] n377 INVx8_ASAP7_75t_R
XU1750 VSS VDD in_data4[30] n376 INVx8_ASAP7_75t_R
XU1751 VSS VDD in_data4[29] n375 INVx8_ASAP7_75t_R
XU1752 VSS VDD in_data4[28] n374 INVx8_ASAP7_75t_R
XU1753 VSS VDD in_data4[27] n373 INVx8_ASAP7_75t_R
XU1754 VSS VDD in_data4[26] n372 INVx8_ASAP7_75t_R
XU1755 VSS VDD in_data4[25] n371 INVx8_ASAP7_75t_R
XU1756 VSS VDD in_data4[24] n370 INVx8_ASAP7_75t_R
XU1757 VSS VDD in_data4[23] n369 INVx8_ASAP7_75t_R
XU1758 VSS VDD in_data4[22] n368 INVx8_ASAP7_75t_R
XU1759 VSS VDD in_data4[21] n367 INVx8_ASAP7_75t_R
XU1760 VSS VDD in_data4[20] n366 INVx8_ASAP7_75t_R
XU1761 VSS VDD in_data4[19] n365 INVx8_ASAP7_75t_R
XU1762 VSS VDD in_data4[18] n364 INVx8_ASAP7_75t_R
XU1763 VSS VDD in_data4[17] n363 INVx8_ASAP7_75t_R
XU1764 VSS VDD in_data4[16] n362 INVx8_ASAP7_75t_R
XU1765 VSS VDD in_data4[15] n361 INVx8_ASAP7_75t_R
XU1766 VSS VDD in_data4[14] n360 INVx8_ASAP7_75t_R
XU1767 VSS VDD in_data4[13] n359 INVx8_ASAP7_75t_R
XU1768 VSS VDD in_data4[12] n358 INVx8_ASAP7_75t_R
XU1769 VSS VDD in_data4[11] n357 INVx8_ASAP7_75t_R
XU1770 VSS VDD in_data4[10] n356 INVx8_ASAP7_75t_R
XU1771 VSS VDD in_data4[9] n355 INVx8_ASAP7_75t_R
XU1772 VSS VDD in_data4[8] n354 INVx8_ASAP7_75t_R
XU1773 VSS VDD in_data4[7] n353 INVx8_ASAP7_75t_R
XU1774 VSS VDD in_data4[6] n352 INVx8_ASAP7_75t_R
XU1775 VSS VDD in_data4[5] n351 INVx8_ASAP7_75t_R
XU1776 VSS VDD in_data4[4] n350 INVx8_ASAP7_75t_R
XU1777 VSS VDD in_data4[3] n349 INVx8_ASAP7_75t_R
XU1778 VSS VDD in_data4[2] n348 INVx8_ASAP7_75t_R
XU1779 VSS VDD in_data4[1] n347 INVx8_ASAP7_75t_R
XU1780 VSS VDD in_data4[0] n346 INVx8_ASAP7_75t_R
XU950 VSS VDD n335 O4[4] INVxp33_ASAP7_75t_R
XU951 VSS VDD n313 O2[8] INVxp33_ASAP7_75t_R
XU952 VSS VDD n339 O4[8] INVxp33_ASAP7_75t_R
XU953 VSS VDD n316 O2[11] INVxp33_ASAP7_75t_R
XU954 VSS VDD n336 O4[5] INVxp33_ASAP7_75t_R
XU955 VSS VDD n340 O4[9] INVxp33_ASAP7_75t_R
XU956 VSS VDD n337 O4[6] INVxp33_ASAP7_75t_R
XU957 VSS VDD n315 O2[10] INVxp33_ASAP7_75t_R
XU958 VSS VDD n338 O4[7] INVxp33_ASAP7_75t_R
XU959 VSS VDD n312 O2[7] INVxp33_ASAP7_75t_R
XU960 VSS VDD n314 O2[9] INVxp33_ASAP7_75t_R
XU961 VSS VDD n311 O2[6] INVxp33_ASAP7_75t_R
XU962 VSS VDD n341 O4[10] INVxp33_ASAP7_75t_R
XU963 VSS VDD n292 O3[0] INVxp33_ASAP7_75t_R
XU964 VSS VDD n293 O3[1] INVxp33_ASAP7_75t_R
XU965 VSS VDD n294 O3[2] INVxp33_ASAP7_75t_R
XU966 VSS VDD n295 O3[3] INVxp33_ASAP7_75t_R
XU967 VSS VDD n322 O1[4] INVxp33_ASAP7_75t_R
XU968 VSS VDD n296 O3[4] INVxp33_ASAP7_75t_R
XU969 VSS VDD n323 O1[5] INVxp33_ASAP7_75t_R
XU970 VSS VDD n324 O1[6] INVxp33_ASAP7_75t_R
XU971 VSS VDD n297 O3[5] INVxp33_ASAP7_75t_R
XU972 VSS VDD n325 O1[7] INVxp33_ASAP7_75t_R
XU973 VSS VDD n326 O1[8] INVxp33_ASAP7_75t_R
XU974 VSS VDD n327 O1[9] INVxp33_ASAP7_75t_R
XU975 VSS VDD n298 O3[6] INVxp33_ASAP7_75t_R
XU976 VSS VDD n328 O1[10] INVxp33_ASAP7_75t_R
XU977 VSS VDD n299 O3[7] INVxp33_ASAP7_75t_R
XU978 VSS VDD n329 O1[11] INVxp33_ASAP7_75t_R
XU979 VSS VDD n300 O3[8] INVxp33_ASAP7_75t_R
XU980 VSS VDD n330 O1[12] INVxp33_ASAP7_75t_R
XU981 VSS VDD n291 out_valid INVxp33_ASAP7_75t_R
XU982 VSS VDD n334 O4[3] INVxp33_ASAP7_75t_R
XU983 VSS VDD n317 O2[12] INVxp33_ASAP7_75t_R
XU984 VSS VDD n333 O4[2] INVxp33_ASAP7_75t_R
XU985 VSS VDD n332 O4[1] INVxp33_ASAP7_75t_R
XU986 VSS VDD n318 O1[0] INVxp33_ASAP7_75t_R
XU987 VSS VDD n331 O4[0] INVxp33_ASAP7_75t_R
XU988 VSS VDD n310 O2[5] INVxp33_ASAP7_75t_R
XU989 VSS VDD n309 O2[4] INVxp33_ASAP7_75t_R
XU990 VSS VDD n308 O2[3] INVxp33_ASAP7_75t_R
XU991 VSS VDD n307 O2[2] INVxp33_ASAP7_75t_R
XU992 VSS VDD n306 O2[1] INVxp33_ASAP7_75t_R
XU993 VSS VDD n305 O2[0] INVxp33_ASAP7_75t_R
XU994 VSS VDD n319 O1[1] INVxp33_ASAP7_75t_R
XU995 VSS VDD n304 O3[12] INVxp33_ASAP7_75t_R
XU996 VSS VDD n303 O3[11] INVxp33_ASAP7_75t_R
XU997 VSS VDD n302 O3[10] INVxp33_ASAP7_75t_R
XU998 VSS VDD n301 O3[9] INVxp33_ASAP7_75t_R
XU999 VSS VDD n320 O1[2] INVxp33_ASAP7_75t_R
XU1000 VSS VDD n342 O4[11] INVxp33_ASAP7_75t_R
XU1001 VSS VDD n321 O1[3] INVxp33_ASAP7_75t_R
XU1002 VSS VDD n343 O4[12] INVxp33_ASAP7_75t_R
XU942 VSS VDD DP_OP_656J1_124_1759_n67 n1309 INVxp67_ASAP7_75t_R
XU943 VSS VDD DP_OP_654J1_122_1759_n67 n1285 INVxp67_ASAP7_75t_R
XU944 VSS VDD DP_OP_655J1_123_1759_n67 n1301 INVxp67_ASAP7_75t_R
XU945 VSS VDD DP_OP_657J1_125_1759_n67 n1293 INVxp67_ASAP7_75t_R
XU1129 VSS VDD DP_OP_654J1_122_1759_n194 n1141 n1002 n910 MAJIxp5_ASAP7_75t_R
XU1130 VSS VDD DP_OP_657J1_125_1759_n194 n1149 n995 n911 MAJIxp5_ASAP7_75t_R
XU1131 VSS VDD DP_OP_656J1_124_1759_n194 n1123 n993 n912 MAJIxp5_ASAP7_75t_R
XU1132 VSS VDD DP_OP_655J1_123_1759_n194 n1132 n1004 n913 MAJIxp5_ASAP7_75t_R
XU1133 VSS VDD DP_OP_655J1_123_1759_n87 DP_OP_655J1_123_1759_n73 n1233 n914 MAJIxp5_ASAP7_75t_R
XU1134 VSS VDD DP_OP_656J1_124_1759_n87 DP_OP_656J1_124_1759_n73 n1241 n915 MAJIxp5_ASAP7_75t_R
XU1135 VSS VDD DP_OP_654J1_122_1759_n87 DP_OP_654J1_122_1759_n73 n1225 n916 MAJIxp5_ASAP7_75t_R
XU1138 VSS VDD DP_OP_657J1_125_1759_n87 DP_OP_657J1_125_1759_n73 n1217 n917 MAJIxp5_ASAP7_75t_R
XU1789 VSS VDD DP_OP_657J1_125_1759_n77 DP_OP_657J1_125_1759_n75 DP_OP_657J1_125_1759_n71 n1053 MAJIxp5_ASAP7_75t_R
XU1790 VSS VDD DP_OP_654J1_122_1759_n77 DP_OP_654J1_122_1759_n75 DP_OP_654J1_122_1759_n71 n1054 MAJIxp5_ASAP7_75t_R
XU1791 VSS VDD DP_OP_655J1_123_1759_n77 DP_OP_655J1_123_1759_n75 DP_OP_655J1_123_1759_n71 n1055 MAJIxp5_ASAP7_75t_R
XU1792 VSS VDD DP_OP_656J1_124_1759_n77 DP_OP_656J1_124_1759_n75 DP_OP_656J1_124_1759_n71 n1056 MAJIxp5_ASAP7_75t_R
XU1839 VSS VDD DP_OP_654J1_122_1759_n308 DP_OP_654J1_122_1759_n306 DP_OP_654J1_122_1759_n310 n1091 MAJIxp5_ASAP7_75t_R
XU1844 VSS VDD DP_OP_655J1_123_1759_n308 DP_OP_655J1_123_1759_n306 DP_OP_655J1_123_1759_n310 n1098 MAJIxp5_ASAP7_75t_R
XU1849 VSS VDD DP_OP_657J1_125_1759_n308 DP_OP_657J1_125_1759_n306 DP_OP_657J1_125_1759_n310 n1112 MAJIxp5_ASAP7_75t_R
XU1854 VSS VDD DP_OP_656J1_124_1759_n308 DP_OP_656J1_124_1759_n306 DP_OP_656J1_124_1759_n310 n1105 MAJIxp5_ASAP7_75t_R
XU1859 VSS VDD n1091 DP_OP_654J1_122_1759_n258 n1019 n1141 MAJIxp5_ASAP7_75t_R
XU1866 VSS VDD n1098 DP_OP_655J1_123_1759_n258 n1021 n1132 MAJIxp5_ASAP7_75t_R
XU1873 VSS VDD n1105 DP_OP_656J1_124_1759_n258 n1023 n1123 MAJIxp5_ASAP7_75t_R
XU1880 VSS VDD n1112 DP_OP_657J1_125_1759_n258 n1016 n1149 MAJIxp5_ASAP7_75t_R
XU1886 VSS VDD n1120 n1121 n1119 n1162 MAJIxp5_ASAP7_75t_R
XU1891 VSS VDD n1129 n1130 n1128 n1169 MAJIxp5_ASAP7_75t_R
XU1897 VSS VDD n1138 n1139 n1137 n1176 MAJIxp5_ASAP7_75t_R
XU1903 VSS VDD n1146 n1147 n956 n1155 MAJIxp5_ASAP7_75t_R
XU1910 VSS VDD DP_OP_657J1_125_1759_n122 DP_OP_657J1_125_1759_n124 n911 n1186 MAJIxp5_ASAP7_75t_R
XU1912 VSS VDD n1155 n1154 n265 n1183 MAJIxp5_ASAP7_75t_R
XU1917 VSS VDD DP_OP_656J1_124_1759_n122 DP_OP_656J1_124_1759_n124 n912 n1203 MAJIxp5_ASAP7_75t_R
XU1919 VSS VDD n1162 n1161 n187 n1200 MAJIxp5_ASAP7_75t_R
XU1924 VSS VDD DP_OP_655J1_123_1759_n122 DP_OP_655J1_123_1759_n124 n913 n1212 MAJIxp5_ASAP7_75t_R
XU1926 VSS VDD n1169 n1168 n213 n1209 MAJIxp5_ASAP7_75t_R
XU1931 VSS VDD DP_OP_654J1_122_1759_n122 DP_OP_654J1_122_1759_n124 n910 n1194 MAJIxp5_ASAP7_75t_R
XU1933 VSS VDD n1176 n1175 n239 n1191 MAJIxp5_ASAP7_75t_R
XU1937 VSS VDD n1183 n1184 n1182 n1219 MAJIxp5_ASAP7_75t_R
XU1942 VSS VDD n1191 n1192 n957 n1227 MAJIxp5_ASAP7_75t_R
XU1947 VSS VDD n1200 n1201 n1199 n1243 MAJIxp5_ASAP7_75t_R
XU1952 VSS VDD n1209 n1210 n1208 n1235 MAJIxp5_ASAP7_75t_R
XU1959 VSS VDD n269 n1218 n1219 n1250 MAJIxp5_ASAP7_75t_R
XU1965 VSS VDD n243 n1226 n1227 n1259 MAJIxp5_ASAP7_75t_R
XU1971 VSS VDD n217 n1234 n1235 n1268 MAJIxp5_ASAP7_75t_R
XU1977 VSS VDD n191 n1242 n1243 n1277 MAJIxp5_ASAP7_75t_R
XU1981 VSS VDD n1250 n1251 n1042 n1296 MAJIxp5_ASAP7_75t_R
XU1984 VSS VDD DP_OP_657J1_125_1759_n72 DP_OP_657J1_125_1759_n68 n1253 n1294 MAJIxp5_ASAP7_75t_R
XU1987 VSS VDD n1259 n1260 n1043 n1288 MAJIxp5_ASAP7_75t_R
XU1990 VSS VDD DP_OP_654J1_122_1759_n72 DP_OP_654J1_122_1759_n68 n1262 n1286 MAJIxp5_ASAP7_75t_R
XU1993 VSS VDD n1268 n1269 n1267 n1304 MAJIxp5_ASAP7_75t_R
XU1996 VSS VDD DP_OP_655J1_123_1759_n72 DP_OP_655J1_123_1759_n68 n1271 n1302 MAJIxp5_ASAP7_75t_R
XU1999 VSS VDD n1277 n1278 n1044 n1312 MAJIxp5_ASAP7_75t_R
XU2002 VSS VDD DP_OP_656J1_124_1759_n72 DP_OP_656J1_124_1759_n68 n1280 n1310 MAJIxp5_ASAP7_75t_R
XU2005 VSS VDD n1286 DP_OP_654J1_122_1759_n70 n1285 n1363 MAJIxp5_ASAP7_75t_R
XU2006 VSS VDD n247 n1287 n1288 n1360 MAJIxp5_ASAP7_75t_R
XU2007 VSS VDD n1363 n1360 n1361 n1289 MAJIxp5_ASAP7_75t_R
XU2011 VSS VDD n1294 DP_OP_657J1_125_1759_n70 n1293 n1355 MAJIxp5_ASAP7_75t_R
XU2012 VSS VDD n273 n1295 n1296 n1352 MAJIxp5_ASAP7_75t_R
XU2013 VSS VDD n1355 n1352 n1353 n1297 MAJIxp5_ASAP7_75t_R
XU2016 VSS VDD n1302 DP_OP_655J1_123_1759_n70 n1301 n1347 MAJIxp5_ASAP7_75t_R
XU2017 VSS VDD n221 n1303 n1304 n1345 MAJIxp5_ASAP7_75t_R
XU2018 VSS VDD n1347 n1345 n955 n1305 MAJIxp5_ASAP7_75t_R
XU2021 VSS VDD n1310 DP_OP_656J1_124_1759_n70 n1309 n1340 MAJIxp5_ASAP7_75t_R
XU2022 VSS VDD n195 n1311 n1312 n1337 MAJIxp5_ASAP7_75t_R
XU2023 VSS VDD n1340 n1337 n1338 n1313 MAJIxp5_ASAP7_75t_R
XU912 VSS VDD n989 n1194 DP_OP_654J1_122_1759_n88 n1225 MAJx2_ASAP7_75t_R
XU913 VSS VDD n997 n1212 DP_OP_655J1_123_1759_n88 n1233 MAJx2_ASAP7_75t_R
XU914 VSS VDD n999 n1186 DP_OP_657J1_125_1759_n88 n1217 MAJx2_ASAP7_75t_R
XU915 VSS VDD n991 n1203 DP_OP_656J1_124_1759_n88 n1241 MAJx2_ASAP7_75t_R
XU1024 VSS VDD n993 DP_OP_656J1_124_1759_n194 n1123 n935 MAJx2_ASAP7_75t_R
XU1025 VSS VDD n1004 DP_OP_655J1_123_1759_n194 n1132 n936 MAJx2_ASAP7_75t_R
XU1026 VSS VDD n1002 DP_OP_654J1_122_1759_n194 n1141 n933 MAJx2_ASAP7_75t_R
XU1027 VSS VDD n995 DP_OP_657J1_125_1759_n194 n1149 n934 MAJx2_ASAP7_75t_R
XU1174 VSS VDD n1217 DP_OP_657J1_125_1759_n87 DP_OP_657J1_125_1759_n73 n1253 MAJx2_ASAP7_75t_R
XU1175 VSS VDD n1225 DP_OP_654J1_122_1759_n87 DP_OP_654J1_122_1759_n73 n1262 MAJx2_ASAP7_75t_R
XU1176 VSS VDD n1233 DP_OP_655J1_123_1759_n87 DP_OP_655J1_123_1759_n73 n1271 MAJx2_ASAP7_75t_R
XU1177 VSS VDD n1241 DP_OP_656J1_124_1759_n87 DP_OP_656J1_124_1759_n73 n1280 MAJx2_ASAP7_75t_R
XU1003 VSS VDD n1344 n1343 n200 NAND2xp33_ASAP7_75t_R
XU1004 VSS VDD n1383 n1382 n206 NAND2xp33_ASAP7_75t_R
XU1005 VSS VDD n203 n1380 n1381 NAND2xp33_ASAP7_75t_R
XU1006 VSS VDD n1351 n1350 n226 NAND2xp33_ASAP7_75t_R
XU1007 VSS VDD n229 n1368 n1369 NAND2xp33_ASAP7_75t_R
XU1008 VSS VDD n1367 n1366 n252 NAND2xp33_ASAP7_75t_R
XU1009 VSS VDD n1375 n1374 n258 NAND2xp33_ASAP7_75t_R
XU1010 VSS VDD n255 n1372 n1373 NAND2xp33_ASAP7_75t_R
XU1011 VSS VDD n1359 n1358 n278 NAND2xp33_ASAP7_75t_R
XU1012 VSS VDD n1379 n1378 n284 NAND2xp33_ASAP7_75t_R
XU1013 VSS VDD n281 n1376 n1377 NAND2xp33_ASAP7_75t_R
XU1014 VSS VDD in_data2_dff[121] in_data2_dff[113] DP_OP_655J1_123_1759_n227 NAND2xp33_ASAP7_75t_R
XU1015 VSS VDD in_data2_dff[122] in_data2_dff[114] DP_OP_655J1_123_1759_n165 NAND2xp33_ASAP7_75t_R
XU1016 VSS VDD in_data1_dff[121] in_data1_dff[113] DP_OP_654J1_122_1759_n227 NAND2xp33_ASAP7_75t_R
XU1017 VSS VDD in_data4_dff[121] in_data4_dff[113] DP_OP_657J1_125_1759_n227 NAND2xp33_ASAP7_75t_R
XU1018 VSS VDD in_data4_dff[122] in_data4_dff[114] DP_OP_657J1_125_1759_n165 NAND2xp33_ASAP7_75t_R
XU1019 VSS VDD in_data3_dff[112] in_data3_dff[104] DP_OP_656J1_124_1759_n279 NAND2xp33_ASAP7_75t_R
XU1020 VSS VDD in_data3_dff[123] in_data3_dff[115] n1403 NAND2xp33_ASAP7_75t_R
XU1021 VSS VDD in_data2_dff[112] in_data2_dff[104] DP_OP_655J1_123_1759_n279 NAND2xp33_ASAP7_75t_R
XU1022 VSS VDD in_data1_dff[123] in_data1_dff[115] n1401 NAND2xp33_ASAP7_75t_R
XU1023 VSS VDD in_data4_dff[112] in_data4_dff[104] DP_OP_657J1_125_1759_n279 NAND2xp33_ASAP7_75t_R
XU1028 VSS VDD n1111 n1110 n188 NAND2xp33_ASAP7_75t_R
XU1029 VSS VDD n1167 n1166 n192 NAND2xp33_ASAP7_75t_R
XU1030 VSS VDD n1248 n1247 n196 NAND2xp33_ASAP7_75t_R
XU1031 VSS VDD n1313 n199 n1314 NAND2xp33_ASAP7_75t_R
XU1032 VSS VDD n1326 n1325 n204 NAND2xp33_ASAP7_75t_R
XU1033 VSS VDD n1387 n1386 n208 NAND2xp33_ASAP7_75t_R
XU1034 VSS VDD n1104 n1103 n214 NAND2xp33_ASAP7_75t_R
XU1035 VSS VDD n1174 n1173 n218 NAND2xp33_ASAP7_75t_R
XU1036 VSS VDD n1240 n1239 n222 NAND2xp33_ASAP7_75t_R
XU1037 VSS VDD n1305 n225 n1306 NAND2xp33_ASAP7_75t_R
XU1038 VSS VDD n1321 n1320 n230 NAND2xp33_ASAP7_75t_R
XU1039 VSS VDD n1391 n1390 n234 NAND2xp33_ASAP7_75t_R
XU1040 VSS VDD n1097 n1096 n240 NAND2xp33_ASAP7_75t_R
XU1041 VSS VDD n1181 n1180 n244 NAND2xp33_ASAP7_75t_R
XU1042 VSS VDD n1232 n1231 n248 NAND2xp33_ASAP7_75t_R
XU1043 VSS VDD n1289 n251 n1290 NAND2xp33_ASAP7_75t_R
XU1044 VSS VDD n1331 n1330 n256 NAND2xp33_ASAP7_75t_R
XU1045 VSS VDD n1395 n1394 n260 NAND2xp33_ASAP7_75t_R
XU1046 VSS VDD n1398 n1393 n1395 NAND2xp33_ASAP7_75t_R
XU1047 VSS VDD n1118 n1117 n266 NAND2xp33_ASAP7_75t_R
XU1048 VSS VDD n1160 n1159 n270 NAND2xp33_ASAP7_75t_R
XU1049 VSS VDD n1224 n1223 n274 NAND2xp33_ASAP7_75t_R
XU1050 VSS VDD n1297 n277 n1298 NAND2xp33_ASAP7_75t_R
XU1051 VSS VDD n1336 n1335 n282 NAND2xp33_ASAP7_75t_R
XU1052 VSS VDD n1400 n1399 n286 NAND2xp33_ASAP7_75t_R
XU1053 VSS VDD n1398 n1397 n1400 NAND2xp33_ASAP7_75t_R
XU1054 VSS VDD n861 n1143 n1145 NAND2xp33_ASAP7_75t_R
XU1055 VSS VDD n861 n1172 n1173 NAND2xp33_ASAP7_75t_R
XU1056 VSS VDD n861 n1088 n1090 NAND2xp33_ASAP7_75t_R
XU1057 VSS VDD n861 n1158 n1159 NAND2xp33_ASAP7_75t_R
XU1058 VSS VDD n289 n287 n984 NAND2xp33_ASAP7_75t_R
XU1060 VSS VDD n861 n1238 n1239 NAND2xp33_ASAP7_75t_R
XU1061 VSS VDD n861 n1342 n1343 NAND2xp33_ASAP7_75t_R
XU1062 VSS VDD n861 n1357 n1358 NAND2xp33_ASAP7_75t_R
XU1063 VSS VDD n860 n1165 n1166 NAND2xp33_ASAP7_75t_R
XU1064 VSS VDD n860 n1230 n1231 NAND2xp33_ASAP7_75t_R
XU1065 VSS VDD n861 n1246 n1247 NAND2xp33_ASAP7_75t_R
XU1066 VSS VDD n860 n1109 n1110 NAND2xp33_ASAP7_75t_R
XU1067 VSS VDD n861 n1102 n1103 NAND2xp33_ASAP7_75t_R
XU1068 VSS VDD n860 n1080 n1082 NAND2xp33_ASAP7_75t_R
XU1069 VSS VDD n861 n1255 n1257 NAND2xp33_ASAP7_75t_R
XU1070 VSS VDD n861 n1264 n1266 NAND2xp33_ASAP7_75t_R
XU1071 VSS VDD n861 n1273 n1275 NAND2xp33_ASAP7_75t_R
XU1072 VSS VDD n860 n1125 n1127 NAND2xp33_ASAP7_75t_R
XU1073 VSS VDD n861 n1151 n1153 NAND2xp33_ASAP7_75t_R
XU1074 VSS VDD n860 n1196 n1198 NAND2xp33_ASAP7_75t_R
XU1075 VSS VDD n861 n1188 n1190 NAND2xp33_ASAP7_75t_R
XU1076 VSS VDD n861 n1214 n1216 NAND2xp33_ASAP7_75t_R
XU1077 VSS VDD n861 n1222 n1223 NAND2xp33_ASAP7_75t_R
XU1078 VSS VDD n860 n1095 n1096 NAND2xp33_ASAP7_75t_R
XU1079 VSS VDD n861 n1076 n1078 NAND2xp33_ASAP7_75t_R
XU1080 VSS VDD n861 n1205 n1207 NAND2xp33_ASAP7_75t_R
XU1158 VSS VDD n1145 n1144 n242 NAND2xp33_ASAP7_75t_R
XU1159 VSS VDD n1292 n1291 n254 NAND2xp33_ASAP7_75t_R
XU1160 VSS VDD n1086 n1085 n264 NAND2xp33_ASAP7_75t_R
XU1161 VSS VDD n1300 n1299 n280 NAND2xp33_ASAP7_75t_R
XU1162 VSS VDD n1257 n1256 n276 NAND2xp33_ASAP7_75t_R
XU1163 VSS VDD n1275 n1274 n224 NAND2xp33_ASAP7_75t_R
XU1164 VSS VDD n1308 n1307 n228 NAND2xp33_ASAP7_75t_R
XU1165 VSS VDD n1266 n1265 n250 NAND2xp33_ASAP7_75t_R
XU1166 VSS VDD n1153 n1152 n268 NAND2xp33_ASAP7_75t_R
XU1167 VSS VDD n1082 n1081 n212 NAND2xp33_ASAP7_75t_R
XU1168 VSS VDD n1136 n1135 n216 NAND2xp33_ASAP7_75t_R
XU1169 VSS VDD n1216 n1215 n220 NAND2xp33_ASAP7_75t_R
XU1170 VSS VDD n1078 n1077 n238 NAND2xp33_ASAP7_75t_R
XU1171 VSS VDD n1090 n1089 n186 NAND2xp33_ASAP7_75t_R
XU1172 VSS VDD n1127 n1126 n190 NAND2xp33_ASAP7_75t_R
XU1173 VSS VDD n1284 n1283 n198 NAND2xp33_ASAP7_75t_R
XU1229 VSS VDD n1207 n1206 n194 NAND2xp33_ASAP7_75t_R
XU1231 VSS VDD n1198 n1197 n246 NAND2xp33_ASAP7_75t_R
XU1233 VSS VDD n1190 n1189 n272 NAND2xp33_ASAP7_75t_R
XU1245 VSS VDD n861 n1365 n1366 NAND2xp33_ASAP7_75t_R
XU1248 VSS VDD n860 n1134 n1136 NAND2xp33_ASAP7_75t_R
XU1249 VSS VDD n860 n1282 n1284 NAND2xp33_ASAP7_75t_R
XU1250 VSS VDD n861 n1116 n1117 NAND2xp33_ASAP7_75t_R
XU1251 VSS VDD n861 n1349 n1350 NAND2xp33_ASAP7_75t_R
XU1252 VSS VDD n861 n1179 n1180 NAND2xp33_ASAP7_75t_R
XU1781 VSS VDD n1045 n1038 n1334 NAND2xp33_ASAP7_75t_R
XU1782 VSS VDD n1046 n1039 n1329 NAND2xp33_ASAP7_75t_R
XU1783 VSS VDD n1047 n1040 n1319 NAND2xp33_ASAP7_75t_R
XU1784 VSS VDD n1048 n1041 n1324 NAND2xp33_ASAP7_75t_R
XU1785 VSS VDD n1332 n1333 n1376 NAND2xp33_ASAP7_75t_R
XU1786 VSS VDD n1327 n1328 n1372 NAND2xp33_ASAP7_75t_R
XU1787 VSS VDD n1317 n1318 n1368 NAND2xp33_ASAP7_75t_R
XU1788 VSS VDD n1322 n1323 n1380 NAND2xp33_ASAP7_75t_R
XU1793 VSS VDD n1338 n1057 n1283 NAND2xp33_ASAP7_75t_R
XU1794 VSS VDD n955 n1057 n1274 NAND2xp33_ASAP7_75t_R
XU1795 VSS VDD n1353 n1057 n1256 NAND2xp33_ASAP7_75t_R
XU1796 VSS VDD n1044 n1057 n1206 NAND2xp33_ASAP7_75t_R
XU1797 VSS VDD n1043 n1057 n1197 NAND2xp33_ASAP7_75t_R
XU1798 VSS VDD n1057 n1042 n1189 NAND2xp33_ASAP7_75t_R
XU1799 VSS VDD n1317 n1057 n1307 NAND2xp33_ASAP7_75t_R
XU1800 VSS VDD n1327 n1057 n1291 NAND2xp33_ASAP7_75t_R
XU1801 VSS VDD n1322 n1057 n1315 NAND2xp33_ASAP7_75t_R
XU1802 VSS VDD in_data3_dff[121] in_data3_dff[113] DP_OP_656J1_124_1759_n227 NAND2xp33_ASAP7_75t_R
XU1803 VSS VDD in_data3_dff[122] in_data3_dff[114] DP_OP_656J1_124_1759_n165 NAND2xp33_ASAP7_75t_R
XU1804 VSS VDD in_data2_dff[123] in_data2_dff[115] n1402 NAND2xp33_ASAP7_75t_R
XU1805 VSS VDD in_data1_dff[112] in_data1_dff[104] DP_OP_654J1_122_1759_n279 NAND2xp33_ASAP7_75t_R
XU1806 VSS VDD in_data1_dff[122] in_data1_dff[114] DP_OP_654J1_122_1759_n165 NAND2xp33_ASAP7_75t_R
XU1807 VSS VDD in_data4_dff[123] in_data4_dff[115] n1404 NAND2xp33_ASAP7_75t_R
XU1808 VSS VDD n860 n1067 n1068 NAND2xp33_ASAP7_75t_R
XU1809 VSS VDD n1199 n1057 n1126 NAND2xp33_ASAP7_75t_R
XU1810 VSS VDD n1398 n1385 n1387 NAND2xp33_ASAP7_75t_R
XU1811 VSS VDD n1267 n1057 n1215 NAND2xp33_ASAP7_75t_R
XU1812 VSS VDD n1398 n1389 n1391 NAND2xp33_ASAP7_75t_R
XU1813 VSS VDD n1057 n1361 n1265 NAND2xp33_ASAP7_75t_R
XU1814 VSS VDD n860 n1084 n1086 NAND2xp33_ASAP7_75t_R
XU1815 VSS VDD n1332 n1057 n1299 NAND2xp33_ASAP7_75t_R
XU1816 VSS VDD n1069 n1068 n184 NAND2xp33_ASAP7_75t_R
XU1817 VSS VDD n1316 n1315 n202 NAND2xp33_ASAP7_75t_R
XU1818 VSS VDD n1371 n1370 n232 NAND2xp33_ASAP7_75t_R
XU1819 VSS VDD n1061 n1060 n262 NAND2xp33_ASAP7_75t_R
XU1824 VSS VDD n861 n1059 n1060 NAND2xp33_ASAP7_75t_R
XU1828 VSS VDD n860 n1063 n1064 NAND2xp33_ASAP7_75t_R
XU1829 VSS VDD n1065 n1064 n210 NAND2xp33_ASAP7_75t_R
XU1836 VSS VDD n861 n1071 n1072 NAND2xp33_ASAP7_75t_R
XU1837 VSS VDD n1073 n1072 n236 NAND2xp33_ASAP7_75t_R
XU1842 VSS VDD n1137 n1057 n1077 NAND2xp33_ASAP7_75t_R
XU1847 VSS VDD n1128 n1057 n1081 NAND2xp33_ASAP7_75t_R
XU1852 VSS VDD n956 n1057 n1085 NAND2xp33_ASAP7_75t_R
XU1857 VSS VDD n1119 n1057 n1089 NAND2xp33_ASAP7_75t_R
XU1896 VSS VDD n1208 n1057 n1135 NAND2xp33_ASAP7_75t_R
XU1902 VSS VDD n1057 n957 n1144 NAND2xp33_ASAP7_75t_R
XU1908 VSS VDD n1057 n1182 n1152 NAND2xp33_ASAP7_75t_R
XU2010 VSS VDD n1290 n1398 n1039 n1292 NAND3xp33_ASAP7_75t_R
XU2015 VSS VDD n1298 n1398 n1038 n1300 NAND3xp33_ASAP7_75t_R
XU2020 VSS VDD n1306 n1398 n1040 n1308 NAND3xp33_ASAP7_75t_R
XU2025 VSS VDD n1314 n1398 n1041 n1316 NAND3xp33_ASAP7_75t_R
XU2026 VSS VDD n1319 n1398 n1368 n1321 NAND3xp33_ASAP7_75t_R
XU2028 VSS VDD n1324 n1398 n1380 n1326 NAND3xp33_ASAP7_75t_R
XU2030 VSS VDD n1329 n1398 n1372 n1331 NAND3xp33_ASAP7_75t_R
XU2032 VSS VDD n1334 n1398 n1376 n1336 NAND3xp33_ASAP7_75t_R
XU2051 VSS VDD n1369 n1398 n1051 n1371 NAND3xp33_ASAP7_75t_R
XU2054 VSS VDD n1373 n1398 n1050 n1375 NAND3xp33_ASAP7_75t_R
XU2057 VSS VDD n1377 n1398 n1049 n1379 NAND3xp33_ASAP7_75t_R
XU2060 VSS VDD n1381 n1398 n1052 n1383 NAND3xp33_ASAP7_75t_R
XU1081 VSS VDD n344 n984 n863 NOR2xp33_ASAP7_75t_R
XU1838 VSS VDD n1074 n235 n1075 NOR2xp33_ASAP7_75t_R
XU1843 VSS VDD n1074 n209 n1079 NOR2xp33_ASAP7_75t_R
XU1848 VSS VDD n1074 n261 n1083 NOR2xp33_ASAP7_75t_R
XU1853 VSS VDD n1074 n182 n1087 NOR2xp33_ASAP7_75t_R
XU1861 VSS VDD n235 n1092 n1139 NOR2xp33_ASAP7_75t_R
XU1863 VSS VDD n1074 n1093 n1094 NOR2xp33_ASAP7_75t_R
XU1868 VSS VDD n209 n1099 n1130 NOR2xp33_ASAP7_75t_R
XU1870 VSS VDD n1074 n1100 n1101 NOR2xp33_ASAP7_75t_R
XU1875 VSS VDD n182 n1106 n1121 NOR2xp33_ASAP7_75t_R
XU1877 VSS VDD n1074 n1107 n1108 NOR2xp33_ASAP7_75t_R
XU1882 VSS VDD n261 n1113 n1147 NOR2xp33_ASAP7_75t_R
XU1884 VSS VDD n1074 n1114 n1115 NOR2xp33_ASAP7_75t_R
XU1888 VSS VDD n1074 n1122 n1124 NOR2xp33_ASAP7_75t_R
XU1893 VSS VDD n1074 n1131 n1133 NOR2xp33_ASAP7_75t_R
XU1899 VSS VDD n1074 n1140 n1142 NOR2xp33_ASAP7_75t_R
XU1905 VSS VDD n1074 n1148 n1150 NOR2xp33_ASAP7_75t_R
XU1914 VSS VDD n1074 n1156 n1157 NOR2xp33_ASAP7_75t_R
XU1921 VSS VDD n1074 n1163 n1164 NOR2xp33_ASAP7_75t_R
XU1928 VSS VDD n1074 n1170 n1171 NOR2xp33_ASAP7_75t_R
XU1935 VSS VDD n1074 n1177 n1178 NOR2xp33_ASAP7_75t_R
XU1939 VSS VDD n1074 n1185 n1187 NOR2xp33_ASAP7_75t_R
XU1944 VSS VDD n1074 n1193 n1195 NOR2xp33_ASAP7_75t_R
XU1949 VSS VDD n1074 n1202 n1204 NOR2xp33_ASAP7_75t_R
XU1954 VSS VDD n1074 n1211 n1213 NOR2xp33_ASAP7_75t_R
XU1961 VSS VDD n1074 n1220 n1221 NOR2xp33_ASAP7_75t_R
XU1967 VSS VDD n1074 n1228 n1229 NOR2xp33_ASAP7_75t_R
XU1973 VSS VDD n1074 n1236 n1237 NOR2xp33_ASAP7_75t_R
XU1979 VSS VDD n1074 n1244 n1245 NOR2xp33_ASAP7_75t_R
XU1983 VSS VDD n1074 n1252 n1254 NOR2xp33_ASAP7_75t_R
XU1989 VSS VDD n1074 n1261 n1263 NOR2xp33_ASAP7_75t_R
XU1995 VSS VDD n1074 n1270 n1272 NOR2xp33_ASAP7_75t_R
XU2001 VSS VDD n1074 n1279 n1281 NOR2xp33_ASAP7_75t_R
XU2008 VSS VDD n1057 n1074 n1398 NOR2xp33_ASAP7_75t_R
XU2009 VSS VDD n251 n1289 n1328 NOR2xp33_ASAP7_75t_R
XU2014 VSS VDD n277 n1297 n1333 NOR2xp33_ASAP7_75t_R
XU2019 VSS VDD n225 n1305 n1318 NOR2xp33_ASAP7_75t_R
XU2024 VSS VDD n199 n1313 n1323 NOR2xp33_ASAP7_75t_R
XU2036 VSS VDD n1074 n1339 n1341 NOR2xp33_ASAP7_75t_R
XU2040 VSS VDD n1074 n1346 n1348 NOR2xp33_ASAP7_75t_R
XU2044 VSS VDD n1074 n1354 n1356 NOR2xp33_ASAP7_75t_R
XU2048 VSS VDD n1074 n1362 n1364 NOR2xp33_ASAP7_75t_R
XU2050 VSS VDD n229 n1368 n1388 NOR2xp33_ASAP7_75t_R
XU2053 VSS VDD n255 n1372 n1392 NOR2xp33_ASAP7_75t_R
XU2056 VSS VDD n281 n1376 n1396 NOR2xp33_ASAP7_75t_R
XU2059 VSS VDD n203 n1380 n1384 NOR2xp33_ASAP7_75t_R
XU2166 VSS VDD DP_OP_654J1_122_1759_n186 n1401 DP_OP_654J1_122_1759_n116 NOR2xp33_ASAP7_75t_R
XU2172 VSS VDD DP_OP_655J1_123_1759_n186 n1402 DP_OP_655J1_123_1759_n116 NOR2xp33_ASAP7_75t_R
XU2178 VSS VDD DP_OP_656J1_124_1759_n186 n1403 DP_OP_656J1_124_1759_n116 NOR2xp33_ASAP7_75t_R
XU2184 VSS VDD DP_OP_657J1_125_1759_n186 n1404 DP_OP_657J1_125_1759_n116 NOR2xp33_ASAP7_75t_R
XU2190 VSS VDD n261 n862 N1602 NOR2xp33_ASAP7_75t_R
XU2191 VSS VDD n1027 n862 N1603 NOR2xp33_ASAP7_75t_R
XU2192 VSS VDD n862 n265 N1604 NOR2xp33_ASAP7_75t_R
XU2193 VSS VDD n1026 n862 N1605 NOR2xp33_ASAP7_75t_R
XU2194 VSS VDD n269 n862 N1606 NOR2xp33_ASAP7_75t_R
XU2195 VSS VDD n1249 n862 N1607 NOR2xp33_ASAP7_75t_R
XU2196 VSS VDD n273 n862 N1608 NOR2xp33_ASAP7_75t_R
XU2197 VSS VDD n1025 n862 N1609 NOR2xp33_ASAP7_75t_R
XU2198 VSS VDD n277 n862 N1610 NOR2xp33_ASAP7_75t_R
XU2199 VSS VDD n1045 n862 N1611 NOR2xp33_ASAP7_75t_R
XU2200 VSS VDD n281 n862 N1612 NOR2xp33_ASAP7_75t_R
XU2201 VSS VDD n862 n283 N1613 NOR2xp33_ASAP7_75t_R
XU2202 VSS VDD n285 n862 N1614 NOR2xp33_ASAP7_75t_R
XU2203 VSS VDD n182 n862 N1589 NOR2xp33_ASAP7_75t_R
XU2204 VSS VDD n1037 n862 N1590 NOR2xp33_ASAP7_75t_R
XU2205 VSS VDD n862 n187 N1591 NOR2xp33_ASAP7_75t_R
XU2206 VSS VDD n1036 n862 N1592 NOR2xp33_ASAP7_75t_R
XU2207 VSS VDD n191 n862 N1593 NOR2xp33_ASAP7_75t_R
XU2208 VSS VDD n1276 n862 N1594 NOR2xp33_ASAP7_75t_R
XU2209 VSS VDD n862 n195 N1595 NOR2xp33_ASAP7_75t_R
XU2210 VSS VDD n1035 n862 N1596 NOR2xp33_ASAP7_75t_R
XU2211 VSS VDD n199 n862 N1597 NOR2xp33_ASAP7_75t_R
XU2212 VSS VDD n1048 n862 N1598 NOR2xp33_ASAP7_75t_R
XU2213 VSS VDD n862 n203 N1599 NOR2xp33_ASAP7_75t_R
XU2214 VSS VDD n205 n862 N1600 NOR2xp33_ASAP7_75t_R
XU2215 VSS VDD n207 n862 N1601 NOR2xp33_ASAP7_75t_R
XU2216 VSS VDD n209 n862 N1576 NOR2xp33_ASAP7_75t_R
XU2217 VSS VDD n1034 n862 N1577 NOR2xp33_ASAP7_75t_R
XU2218 VSS VDD n213 n862 N1578 NOR2xp33_ASAP7_75t_R
XU2219 VSS VDD n1033 n862 N1579 NOR2xp33_ASAP7_75t_R
XU2220 VSS VDD n217 n862 N1580 NOR2xp33_ASAP7_75t_R
XU2221 VSS VDD n1032 n862 N1581 NOR2xp33_ASAP7_75t_R
XU2222 VSS VDD n221 n862 N1582 NOR2xp33_ASAP7_75t_R
XU2223 VSS VDD n1031 n862 N1583 NOR2xp33_ASAP7_75t_R
XU2224 VSS VDD n225 n862 N1584 NOR2xp33_ASAP7_75t_R
XU2225 VSS VDD n1047 n862 N1585 NOR2xp33_ASAP7_75t_R
XU2226 VSS VDD n229 n862 N1586 NOR2xp33_ASAP7_75t_R
XU2227 VSS VDD n231 n862 N1587 NOR2xp33_ASAP7_75t_R
XU2228 VSS VDD n233 n862 N1588 NOR2xp33_ASAP7_75t_R
XU2229 VSS VDD n235 n862 N1563 NOR2xp33_ASAP7_75t_R
XU2230 VSS VDD n1030 n862 N1564 NOR2xp33_ASAP7_75t_R
XU2231 VSS VDD n862 n239 N1565 NOR2xp33_ASAP7_75t_R
XU2232 VSS VDD n1029 n862 N1566 NOR2xp33_ASAP7_75t_R
XU2233 VSS VDD n862 n243 N1567 NOR2xp33_ASAP7_75t_R
XU2234 VSS VDD n1258 n862 N1568 NOR2xp33_ASAP7_75t_R
XU2235 VSS VDD n247 n862 N1569 NOR2xp33_ASAP7_75t_R
XU2236 VSS VDD n1028 n862 N1570 NOR2xp33_ASAP7_75t_R
XU2237 VSS VDD n251 n862 N1571 NOR2xp33_ASAP7_75t_R
XU2238 VSS VDD n1046 n862 N1572 NOR2xp33_ASAP7_75t_R
XU2239 VSS VDD n255 n862 N1573 NOR2xp33_ASAP7_75t_R
XU2240 VSS VDD n257 n862 N1574 NOR2xp33_ASAP7_75t_R
XU2241 VSS VDD n259 n862 N1575 NOR2xp33_ASAP7_75t_R
XU2243 VSS VDD n1057 n289 n1405 NOR2xp33_ASAP7_75t_R
XU1059 VSS VDD n984 n344 n862 OR2x2_ASAP7_75t_R
XU1178 VSS VDD n1297 n277 n1038 OR2x2_ASAP7_75t_R
XU1179 VSS VDD n1289 n251 n1039 OR2x2_ASAP7_75t_R
XU1180 VSS VDD n1305 n225 n1040 OR2x2_ASAP7_75t_R
XU1181 VSS VDD n1313 n199 n1041 OR2x2_ASAP7_75t_R
XU1182 VSS VDD n1376 n281 n1049 OR2x2_ASAP7_75t_R
XU1183 VSS VDD n1372 n255 n1050 OR2x2_ASAP7_75t_R
XU1184 VSS VDD n1368 n229 n1051 OR2x2_ASAP7_75t_R
XU1185 VSS VDD n1380 n203 n1052 OR2x2_ASAP7_75t_R
XU1821 VSS VDD n261 n861 n1061 OR2x2_ASAP7_75t_R
XU1825 VSS VDD n209 n861 n1065 OR2x2_ASAP7_75t_R
XU1830 VSS VDD n182 n860 n1069 OR2x2_ASAP7_75t_R
XU1833 VSS VDD n235 n861 n1073 OR2x2_ASAP7_75t_R
XU1858 VSS VDD n239 n861 n1097 OR2x2_ASAP7_75t_R
XU1865 VSS VDD n213 n861 n1104 OR2x2_ASAP7_75t_R
XU1872 VSS VDD n187 n860 n1111 OR2x2_ASAP7_75t_R
XU1879 VSS VDD n265 n861 n1118 OR2x2_ASAP7_75t_R
XU1909 VSS VDD n269 n861 n1160 OR2x2_ASAP7_75t_R
XU1916 VSS VDD n191 n861 n1167 OR2x2_ASAP7_75t_R
XU1923 VSS VDD n217 n860 n1174 OR2x2_ASAP7_75t_R
XU1930 VSS VDD n243 n861 n1181 OR2x2_ASAP7_75t_R
XU1957 VSS VDD n273 n861 n1224 OR2x2_ASAP7_75t_R
XU1963 VSS VDD n247 n860 n1232 OR2x2_ASAP7_75t_R
XU1969 VSS VDD n221 n861 n1240 OR2x2_ASAP7_75t_R
XU1975 VSS VDD n195 n861 n1248 OR2x2_ASAP7_75t_R
XU2027 VSS VDD n229 n860 n1320 OR2x2_ASAP7_75t_R
XU2029 VSS VDD n203 n861 n1325 OR2x2_ASAP7_75t_R
XU2031 VSS VDD n255 n860 n1330 OR2x2_ASAP7_75t_R
XU2033 VSS VDD n281 n861 n1335 OR2x2_ASAP7_75t_R
XU2034 VSS VDD n199 n861 n1344 OR2x2_ASAP7_75t_R
XU2038 VSS VDD n225 n861 n1351 OR2x2_ASAP7_75t_R
XU2042 VSS VDD n277 n860 n1359 OR2x2_ASAP7_75t_R
XU2046 VSS VDD n251 n861 n1367 OR2x2_ASAP7_75t_R
XU2052 VSS VDD n231 n861 n1370 OR2x2_ASAP7_75t_R
XU2055 VSS VDD n257 n860 n1374 OR2x2_ASAP7_75t_R
XU2058 VSS VDD n283 n861 n1378 OR2x2_ASAP7_75t_R
XU2061 VSS VDD n205 n860 n1382 OR2x2_ASAP7_75t_R
XU2063 VSS VDD n207 n860 n1386 OR2x2_ASAP7_75t_R
XU2089 VSS VDD n233 n861 n1390 OR2x2_ASAP7_75t_R
XU2115 VSS VDD n259 n860 n1394 OR2x2_ASAP7_75t_R
XU2141 VSS VDD n285 n861 n1399 OR2x2_ASAP7_75t_R
XU1820 VSS VDD n183 TIELOx1_ASAP7_75t_R
XU1822 VSS VDD DP_OP_657J1_125_1759_n310 DP_OP_657J1_125_1759_n308 n1058 XOR2xp5_ASAP7_75t_R
XU1823 VSS VDD DP_OP_657J1_125_1759_n306 n1058 n1059 XOR2xp5_ASAP7_75t_R
XU1826 VSS VDD DP_OP_655J1_123_1759_n310 DP_OP_655J1_123_1759_n308 n1062 XOR2xp5_ASAP7_75t_R
XU1827 VSS VDD DP_OP_655J1_123_1759_n306 n1062 n1063 XOR2xp5_ASAP7_75t_R
XU1831 VSS VDD DP_OP_656J1_124_1759_n310 DP_OP_656J1_124_1759_n308 n1066 XOR2xp5_ASAP7_75t_R
XU1832 VSS VDD DP_OP_656J1_124_1759_n306 n1066 n1067 XOR2xp5_ASAP7_75t_R
XU1834 VSS VDD DP_OP_654J1_122_1759_n310 DP_OP_654J1_122_1759_n308 n1070 XOR2xp5_ASAP7_75t_R
XU1835 VSS VDD DP_OP_654J1_122_1759_n306 n1070 n1071 XOR2xp5_ASAP7_75t_R
XU1864 VSS VDD n1138 n1094 n1095 XOR2xp5_ASAP7_75t_R
XU1871 VSS VDD n1129 n1101 n1102 XOR2xp5_ASAP7_75t_R
XU1878 VSS VDD n1120 n1108 n1109 XOR2xp5_ASAP7_75t_R
XU1885 VSS VDD n1146 n1115 n1116 XOR2xp5_ASAP7_75t_R
XU1915 VSS VDD n1184 n1157 n1158 XOR2xp5_ASAP7_75t_R
XU1922 VSS VDD n1201 n1164 n1165 XOR2xp5_ASAP7_75t_R
XU1929 VSS VDD n1210 n1171 n1172 XOR2xp5_ASAP7_75t_R
XU1936 VSS VDD n1192 n1178 n1179 XOR2xp5_ASAP7_75t_R
XU1962 VSS VDD n1251 n1221 n1222 XOR2xp5_ASAP7_75t_R
XU1968 VSS VDD n1260 n1229 n1230 XOR2xp5_ASAP7_75t_R
XU1974 VSS VDD n1269 n1237 n1238 XOR2xp5_ASAP7_75t_R
XU1980 VSS VDD n1278 n1245 n1246 XOR2xp5_ASAP7_75t_R
XU2037 VSS VDD n1341 n1340 n1342 XOR2xp5_ASAP7_75t_R
XU2041 VSS VDD n1348 n1347 n1349 XOR2xp5_ASAP7_75t_R
XU2045 VSS VDD n1356 n1355 n1357 XOR2xp5_ASAP7_75t_R
XU2049 VSS VDD n1364 n1363 n1365 XOR2xp5_ASAP7_75t_R
XU2167 VSS VDD DP_OP_654J1_122_1759_n186 n1401 DP_OP_654J1_122_1759_n117 XOR2xp5_ASAP7_75t_R
XU2173 VSS VDD DP_OP_655J1_123_1759_n186 n1402 DP_OP_655J1_123_1759_n117 XOR2xp5_ASAP7_75t_R
XU2179 VSS VDD DP_OP_656J1_124_1759_n186 n1403 DP_OP_656J1_124_1759_n117 XOR2xp5_ASAP7_75t_R
XU2185 VSS VDD DP_OP_657J1_125_1759_n186 n1404 DP_OP_657J1_125_1759_n117 XOR2xp5_ASAP7_75t_R
.ENDS
